//: version "1.8.7"

module UC();
//: interface  /sz:(101, 231) /bd:[ Bi0>Op[5:0](34/101) Bi1>Funct[5:0](61/101) Ro0<Branch(32/231) Ro1<Jump(17/231) Ro2<MemRead(50/231) Ro3<MemToRed(66/231) Ro4<ALUCtrl[3:0](174/231) Ro5<MemWrite(85/231) Ro6<ALUSrc(101/231) Ro7<RegWrite(120/231) Ro8<RegDst(209/231) ]
//: enddecls


endmodule

module Mem(MemRead, MemWrite, WriteData, ReadData, Address);
//: interface  /sz:(147, 210) /bd:[ Ti0>MemWrite(86/147) Li0>Adress[31:0](72/210) Li1>WriteData[31:0](148/210) Bi0>MemRead(80/147) Ro0<ReadData[31:0](78/210) ]
output [31:0] ReadData;    //: /sn:0 /dp:1 {0}(596,161)(660,161){1}
//: {2}(664,161)(854,161){3}
//: {4}(662,163)(662,172){5}
supply0 w0;    //: /sn:0 {0}(572,208)(572,188){1}
input [31:0] WriteData;    //: /sn:0 {0}(740,179)(750,179)(750,194)(662,194)(662,188){1}
input MemWrite;    //: /sn:0 {0}(562,71)(579,71)(579,93){1}
//: {2}(581,95)(636,95)(636,180)(657,180){3}
//: {4}(579,97)(579,138){5}
input MemRead;    //: /sn:0 {0}(529,226)(586,226)(586,188){1}
input [31:0] Address;    //: /sn:0 /dp:1 {0}(561,163)(539,163)(539,130)(334,130){1}
//: enddecls

  //: supply0 g4 (w0) @(572,214) /sn:0 /w:[ 0 ]
  //: joint g8 (ReadData) @(662, 161) /w:[ 2 -1 1 4 ]
  //: input g3 (MemRead) @(527,226) /sn:0 /w:[ 0 ]
  //: input g2 (MemWrite) @(560,71) /sn:0 /w:[ 0 ]
  ram g1 (.A(Address), .D(ReadData), .WE(!MemWrite), .OE(!MemRead), .CS(w0));   //: @(579,162) /sn:0 /w:[ 0 0 5 1 1 ]
  //: joint g10 (MemWrite) @(579, 95) /w:[ 2 1 -1 4 ]
  bufif1 g6 (.Z(ReadData), .I(WriteData), .E(MemWrite));   //: @(662,182) /sn:0 /R:1 /w:[ 5 1 3 ]
  //: input g7 (WriteData) @(738,179) /sn:0 /w:[ 0 ]
  //: output g9 (ReadData) @(851,161) /sn:0 /w:[ 3 ]
  //: comment g5 /dolink:0 /link:"" @(370,188) /sn:0
  //: /line:"Negate to write on low cycle"
  //: /end
  //: input g0 (Address) @(332,130) /sn:0 /w:[ 1 ]

endmodule

module fetch(Clk, PCNew, Reset, PCNext, Inst);
//: interface  /sz:(88, 222) /bd:[ Li0>PCNew[31:0](13/222) Li1>Clk(160/222) Li2>Reset(44/222) Ro0<Inst[31:0](159/222) Ro1<PCNext[31:0](38/222) ]
input Clk;    //: /sn:0 {0}(122,387)(184,387)(184,357){1}
input [31:0] PCNew;    //: /sn:0 {0}(124,319)(173,319){1}
output [31:0] Inst;    //: /sn:0 /dp:1 {0}(330,317)(369,317){1}
output [31:0] PCNext;    //: /sn:0 {0}(416,153)(360,153){1}
input Reset;    //: /sn:0 {0}(124,265)(179,265)(179,281){1}
supply0 [31:0] w11;    //: /sn:0 {0}(331,169)(323,169){1}
//: {2}(322,169)(314,169)(314,178){3}
wire Cout;    //: /sn:0 {0}(345,177)(345,187){1}
wire w2;    //: /sn:0 {0}(189,281)(189,153)(212,153){1}
//: {2}(216,153)(323,153)(323,164){3}
//: {4}(214,151)(214,116)(345,116)(345,129){5}
//: {6}(214,155)(214,358)(313,358)(313,344){7}
wire [31:0] x;    //: /sn:0 /dp:4 {0}(194,319)(243,319){1}
//: {2}(247,319)(295,319){3}
//: {4}(245,317)(245,137)(331,137){5}
//: enddecls

  //: input g8 (Clk) @(120,387) /sn:0 /w:[ 0 ]
  //: supply0 g3 (w11) @(314,184) /sn:0 /w:[ 3 ]
  add g2 (.A(w11), .B(x), .S(PCNext), .CI(!w2), .CO(Cout));   //: @(347,153) /sn:0 /R:1 /w:[ 0 5 1 5 0 ]
  register g1 (.Q(x), .D(PCNew), .EN(w2), .CLR(!Reset), .CK(!Clk));   //: @(184,319) /sn:0 /R:1 /w:[ 0 1 0 1 1 ]
  tran g10(.Z(w2), .I(w11[0]));   //: @(323,167) /sn:0 /R:1 /w:[ 3 2 1 ] /ss:0
  //: input g6 (PCNew) @(122,319) /sn:0 /w:[ 0 ]
  //: input g9 (Reset) @(122,265) /sn:0 /w:[ 0 ]
  //: output g7 (PCNext) @(413,153) /sn:0 /w:[ 0 ]
  //: output g12 (Inst) @(366,317) /sn:0 /w:[ 1 ]
  //: joint g5 (x) @(245, 319) /w:[ 2 4 1 -1 ]
  //: joint g11 (w2) @(214, 153) /w:[ 2 4 1 6 ]
  rom g0 (.A(x), .D(Inst), .OE(w2));   //: @(313,318) /sn:0 /w:[ 3 0 7 ] /mem:"/home/milax/Documents/EC/EC_Prac2_V2/mult.mem"

endmodule

module ALU(B, ALUResult, ALUOperation, Zero, A);
//: interface  /sz:(96, 97) /bd:[ Ti0>ALUOperation[3:0](44/96) Li0>B[31:0](65/97) Li1>A[31:0](28/97) Ro0<Zero(20/97) Ro1<ALUResult[31:0](45/97) ]
input [31:0] B;    //: /sn:0 {0}(304,108)(191,108){1}
//: {2}(189,106)(189,90){3}
//: {4}(189,110)(189,171){5}
//: {6}(191,173)(305,173){7}
//: {8}(189,175)(189,273)(212,273){9}
output Zero;    //: /sn:0 {0}(656,238)(628,238){1}
supply0 [30:0] Massa;    //: /sn:0 /dp:1 {0}(406,297)(400,297)(400,284)(376,284){1}
input [31:0] A;    //: /sn:0 /dp:1 {0}(305,168)(167,168){1}
//: {2}(165,166)(165,105){3}
//: {4}(167,103)(304,103){5}
//: {6}(165,101)(165,90){7}
//: {8}(165,170)(165,239)(252,239){9}
input [3:0] ALUOperation;    //: /sn:0 {0}(484,89)(484,161){1}
//: {2}(484,162)(484,197){3}
//: {4}(484,198)(484,207){5}
output [31:0] ALUResult;    //: /sn:0 {0}(656,284)(590,284){1}
//: {2}(588,282)(588,238)(607,238){3}
//: {4}(586,284)(554,284){5}
wire [31:0] AsubB;    //: {0}(281,255)(356,255){1}
//: {2}(357,255)(421,255)(421,290)(525,290){3}
wire [31:0] NotBifSub;    //: /sn:0 {0}(233,271)(252,271){1}
wire neg;    //: /sn:0 /dp:1 {0}(357,259)(357,307)(406,307){1}
wire [31:0] AsltB;    //: {0}(412,302)(525,302){1}
wire sub;    //: /dp:1 {0}(479,198)(268,198){1}
//: {2}(264,198)(202,198)(202,268)(212,268){3}
//: {4}(266,200)(266,231){5}
wire [31:0] AorB;    //: {0}(326,171)(432,171)(432,278)(525,278){1}
wire [1:0] Selector;    //: /dp:1 {0}(488,162)(541,162)(541,261){1}
wire [31:0] AandB;    //: {0}(325,106)(441,106)(441,266)(525,266){1}
wire Overflow;    //: /sn:0 {0}(266,279)(266,309)(307,309){1}
//: enddecls

  //: joint g8 (B) @(189, 108) /w:[ 1 2 -1 4 ]
  and g4 (.I0(A), .I1(B), .Z(AandB));   //: @(315,106) /sn:0 /w:[ 5 0 0 ]
  tran g3(.Z(Selector), .I(ALUOperation[1:0]));   //: @(482,162) /sn:0 /R:2 /w:[ 0 2 1 ] /ss:1
  or OR (.I0(A), .I1(B), .Z(AorB));   //: @(316,171) /sn:0 /w:[ 0 7 0 ]
  //: joint g16 (B) @(189, 173) /w:[ 6 5 -1 8 ]
  add g2 (.A(NotBifSub), .B(A), .S(AsubB), .CI(sub), .CO(Overflow));   //: @(268,255) /sn:0 /R:1 /w:[ 1 9 0 5 0 ]
  //: input g1 (B) @(189,88) /sn:0 /R:3 /w:[ 3 ]
  //: output g18 (ALUResult) @(653,284) /sn:0 /w:[ 0 ]
  //: joint g10 (A) @(165, 103) /w:[ 4 6 -1 3 ]
  mux g6 (.I0(AandB), .I1(AorB), .I2(AsubB), .I3(AsltB), .S(Selector), .Z(ALUResult));   //: @(541,284) /sn:0 /R:1 /w:[ 1 1 3 1 1 5 ] /ss:1 /do:1
  //: joint g7 (A) @(165, 168) /w:[ 1 2 -1 8 ]
  //: input g9 (ALUOperation) @(484,87) /sn:0 /R:3 /w:[ 0 ]
  //: supply0 g12 (Massa) @(370,284) /sn:0 /R:3 /w:[ 1 ]
  tran g11(.Z(sub), .I(ALUOperation[2]));   //: @(482,198) /sn:0 /R:2 /w:[ 0 4 3 ] /ss:0
  tran g14(.Z(neg), .I(AsubB[31]));   //: @(357,253) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  xor g5 (.I0(sub), .I1(B), .Z(NotBifSub));   //: @(223,271) /sn:0 /w:[ 3 9 0 ]
  nor g19 (.I0(ALUResult), .Z(Zero));   //: @(618,238) /sn:0 /w:[ 3 1 ]
  //: output g21 (Zero) @(653,238) /sn:0 /w:[ 0 ]
  //: joint g20 (ALUResult) @(588, 284) /w:[ 1 2 4 -1 ]
  //: input g0 (A) @(165,88) /sn:0 /R:3 /w:[ 7 ]
  //: joint g15 (sub) @(266, 198) /w:[ 1 -1 2 4 ]
  concat g13 (.I0(neg), .I1(Massa), .Z(AsltB));   //: @(411,302) /sn:0 /w:[ 1 0 0 ] /dr:0

endmodule

module EXE(PCNext, ALUResult, Zero, rt, rs, Inm32, BranchTarget, ALUOperation, ALUSrc);
//: interface  /sz:(142, 213) /bd:[ Ti0>ALUOperation[3:0](99/142) Ti1>ALUSrc(36/142) Li0>rt[31:0](114/213) Li1>rs[31:0](81/213) Li2>Inm32[31:0](148/213) Li3>PCNext[31:0](25/213) Ro0<ALUResult[31:0](139/213) Ro1<Zero(57/213) ]
output Zero;    //: /sn:0 {0}(473,294)(333,294){1}
input [31:0] Inm32;    //: /sn:0 {0}(99,165)(119,165){1}
//: {2}(123,165)(283,165){3}
//: {4}(121,167)(121,335)(152,335){5}
input [3:0] ALUOperation;    //: /sn:0 /dp:1 {0}(280,273)(280,230)(96,230){1}
input [31:0] rt;    //: /sn:0 {0}(99,355)(152,355){1}
input ALUSrc;    //: /sn:0 {0}(98,389)(168,389)(168,368){1}
output [31:0] ALUResult;    //: /sn:0 {0}(333,319)(474,319){1}
input [31:0] PCNext;    //: /sn:0 {0}(101,133)(283,133){1}
supply0 CarryIn;    //: /sn:0 /dp:1 {0}(244,85)(297,85)(297,125){1}
output [31:0] BranchTarget;    //: /sn:0 {0}(405,149)(312,149){1}
input [31:0] rs;    //: /sn:0 {0}(98,302)(235,302){1}
wire [31:0] w4;    //: /sn:0 /dp:1 {0}(181,345)(235,345){1}
wire Overflow;    //: /sn:0 /dp:1 {0}(297,173)(297,199)(351,199){1}
//: enddecls

  //: input g8 (PCNext) @(99,133) /sn:0 /w:[ 0 ]
  //: output g4 (ALUResult) @(471,319) /sn:0 /w:[ 1 ]
  //: output g3 (Zero) @(470,294) /sn:0 /w:[ 0 ]
  //: input g2 (rt) @(97,355) /sn:0 /w:[ 0 ]
  //: input g1 (rs) @(96,302) /sn:0 /w:[ 0 ]
  //: supply0 g10 (CarryIn) @(238,85) /sn:0 /R:3 /w:[ 0 ]
  add g6 (.A(Inm32), .B(PCNext), .S(BranchTarget), .CI(CarryIn), .CO(Overflow));   //: @(299,149) /sn:0 /R:1 /w:[ 3 1 1 1 0 ]
  //: input g7 (Inm32) @(97,165) /sn:0 /w:[ 0 ]
  //: output g9 (BranchTarget) @(402,149) /sn:0 /w:[ 0 ]
  //: joint g12 (Inm32) @(121, 165) /w:[ 2 -1 1 4 ]
  mux g11 (.I0(rt), .I1(Inm32), .S(ALUSrc), .Z(w4));   //: @(168,345) /sn:0 /R:1 /w:[ 1 5 1 0 ] /ss:0 /do:0
  //: input g5 (ALUOperation) @(94,230) /sn:0 /w:[ 1 ]
  ALU g0 (.ALUOperation(ALUOperation), .B(w4), .A(rs), .Zero(Zero), .ALUResult(ALUResult));   //: @(236, 274) /sz:(96, 97) /sn:0 /p:[ Ti0>0 Li0>1 Li1>1 Ro0<1 Ro1<0 ]
  //: input g13 (ALUSrc) @(96,389) /sn:0 /w:[ 0 ]

endmodule

module BRegs32x32(Read2, Write, Read1, Data2, Data1, clr, clk, RegWrite, WriteData);
//: interface  /sz:(147, 182) /bd:[ Ti0>clr(66/147) Ti1>clr(66/147) Ti2>clr(66/147) Ti3>clr(66/147) Ti4>clr(66/147) Ti5>clr(66/147) Ti6>clr(66/147) Ti7>clr(66/147) Ti8>clr(66/147) Li0>WriteData[31:0](148/182) Li1>Write[4:0](108/182) Li2>Read2[4:0](72/182) Li3>Read1[4:0](32/182) Li4>Read1[4:0](32/182) Li5>Read2[4:0](72/182) Li6>Write[4:0](108/182) Li7>WriteData[31:0](148/182) Li8>WriteData[31:0](148/182) Li9>Write[4:0](108/182) Li10>Read2[4:0](72/182) Li11>Read1[4:0](32/182) Li12>WriteData[31:0](148/182) Li13>Write[4:0](108/182) Li14>Read2[4:0](72/182) Li15>Read1[4:0](32/182) Li16>Read1[4:0](32/182) Li17>Read2[4:0](72/182) Li18>Write[4:0](108/182) Li19>WriteData[31:0](148/182) Li20>WriteData[31:0](148/182) Li21>Write[4:0](108/182) Li22>Read2[4:0](72/182) Li23>Read1[4:0](32/182) Li24>WriteData[31:0](148/182) Li25>Write[4:0](108/182) Li26>Read2[4:0](72/182) Li27>Read1[4:0](32/182) Li28>Read1[4:0](32/182) Li29>Read2[4:0](72/182) Li30>Write[4:0](108/182) Li31>WriteData[31:0](148/182) Li32>WriteData[31:0](148/182) Li33>Write[4:0](108/182) Li34>Read2[4:0](72/182) Li35>Read1[4:0](32/182) Bi0>RegWrite(40/147) Bi1>clk(108/147) Bi2>clk(108/147) Bi3>RegWrite(40/147) Bi4>RegWrite(40/147) Bi5>clk(108/147) Bi6>RegWrite(40/147) Bi7>clk(108/147) Bi8>clk(108/147) Bi9>RegWrite(40/147) Bi10>RegWrite(40/147) Bi11>clk(108/147) Bi12>RegWrite(40/147) Bi13>clk(108/147) Bi14>clk(108/147) Bi15>RegWrite(40/147) Bi16>RegWrite(40/147) Bi17>clk(108/147) Ro0<Data2[31:0](139/182) Ro1<Data1[31:0](47/182) Ro2<Data1[31:0](47/182) Ro3<Data2[31:0](139/182) Ro4<Data2[31:0](139/182) Ro5<Data1[31:0](47/182) Ro6<Data2[31:0](139/182) Ro7<Data1[31:0](47/182) Ro8<Data1[31:0](47/182) Ro9<Data2[31:0](139/182) Ro10<Data2[31:0](139/182) Ro11<Data1[31:0](47/182) Ro12<Data2[31:0](139/182) Ro13<Data1[31:0](47/182) Ro14<Data1[31:0](47/182) Ro15<Data2[31:0](139/182) Ro16<Data2[31:0](139/182) Ro17<Data1[31:0](47/182) ]
output [31:0] Data2;    //: /sn:0 {0}(668,485)(668,472)(669,472)(669,445){1}
input [4:0] Write;    //: /sn:0 {0}(-238,-38)(-138,-38)(-138,-37)(-66,-37){1}
//: {2}(-65,-37)(-28,-37){3}
//: {4}(-27,-37)(-16,-37){5}
input [31:0] WriteData;    //: /sn:0 {0}(669,157)(669,75)(481,75){1}
//: {2}(477,75)(292,75){3}
//: {4}(288,75)(89,75){5}
//: {6}(85,75)(-104,75)(-104,73)(-237,73){7}
//: {8}(87,77)(87,157){9}
//: {10}(290,77)(290,107)(291,107)(291,152){11}
//: {12}(479,77)(479,157){13}
supply1 w21;    //: /sn:0 {0}(82,3)(57,3)(57,-11){1}
output [31:0] Data1;    //: /sn:0 {0}(59,382)(59,465){1}
input RegWrite;    //: /sn:0 {0}(-237,263)(-71,263){1}
//: {2}(-67,263)(171,263){3}
//: {4}(175,263)(370,263){5}
//: {6}(374,263)(552,263)(552,219)(556,219){7}
//: {8}(372,261)(372,219)(383,219){9}
//: {10}(173,261)(173,214)(183,214){11}
//: {12}(-69,261)(-69,219)(-38,219){13}
input clr;    //: /sn:0 {0}(721,193)(731,193)(731,-83)(543,-83){1}
//: {2}(539,-83)(355,-83){3}
//: {4}(351,-83)(150,-83){5}
//: {6}(146,-83)(-44,-83)(-44,-92)(-235,-92){7}
//: {8}(148,-81)(148,193)(139,193){9}
//: {10}(353,-81)(353,188)(343,188){11}
//: {12}(541,-81)(541,193)(531,193){13}
input clk;    //: /sn:0 {0}(556,214)(542,214)(542,285)(364,285){1}
//: {2}(362,283)(362,214)(383,214){3}
//: {4}(360,285)(167,285){5}
//: {6}(165,283)(165,209)(183,209){7}
//: {8}(163,285)(-56,285){9}
//: {10}(-58,283)(-58,214)(-38,214){11}
//: {12}(-60,285)(-237,285){13}
input [4:0] Read1;    //: {0}(-237,96)(-208,96)(-208,95)(-124,95){1}
//: {2}(-123,95)(-96,95){3}
//: {4}(-95,95)(-78,95){5}
input [4:0] Read2;    //: {0}(-237,145)(-141,145){1}
//: {2}(-140,145)(-123,145)(-123,144)(-94,144){3}
//: {4}(-93,144)(-79,144){5}
wire w16;    //: /sn:0 {0}(39,205)(-50,205)(-50,39)(88,39)(88,19){1}
wire [1:0] w6;    //: /sn:0 {0}(36,369)(-123,369)(-123,99){1}
wire w4;    //: /sn:0 {0}(112,19)(112,46)(370,46)(370,205)(431,205){1}
wire w22;    //: /sn:0 {0}(404,217)(431,217){1}
wire [31:0] w0;    //: /sn:0 {0}(651,416)(651,398)(105,398)(105,228){1}
wire [31:0] R2;    //: {0}(65,353)(65,319)(469,319)(469,228){1}
wire [31:0] w3;    //: /sn:0 {0}(77,353)(77,334)(659,334)(659,228){1}
wire w20;    //: /sn:0 {0}(124,19)(124,29)(556,29)(556,205)(621,205){1}
wire [2:0] w18;    //: /sn:0 {0}(431,180)(402,180)(402,125){1}
//: {2}(404,123)(589,123)(589,180)(621,180){3}
//: {4}(400,123)(279,123)(279,122)(212,122){5}
//: {6}(208,122)(8,122){7}
//: {8}(4,122)(-93,122)(-93,139){9}
//: {10}(6,124)(6,180)(39,180){11}
//: {12}(210,124)(210,175)(243,175){13}
wire [2:0] w19;    //: /sn:0 {0}(431,169)(419,169)(419,109){1}
//: {2}(421,107)(606,107)(606,169)(621,169){3}
//: {4}(417,107)(297,107)(297,106)(231,106){5}
//: {6}(227,106)(25,106){7}
//: {8}(21,106)(-95,106)(-95,99){9}
//: {10}(23,108)(23,169)(39,169){11}
//: {12}(229,108)(229,164)(243,164){13}
wire [1:0] w10;    //: /sn:0 {0}(-140,149)(-140,432)(646,432){1}
wire w23;    //: /sn:0 {0}(577,217)(621,217){1}
wire [2:0] w24;    //: /sn:0 {0}(431,193)(381,193)(381,141){1}
//: {2}(383,139)(568,139)(568,193)(621,193){3}
//: {4}(379,139)(260,139)(260,138)(195,138){5}
//: {6}(191,138)(-13,138){7}
//: {8}(-17,138)(-65,138)(-65,-33){9}
//: {10}(-15,140)(-15,193)(39,193){11}
//: {12}(193,140)(193,188)(243,188){13}
wire w1;    //: /sn:0 {0}(-17,217)(39,217){1}
wire w31;    //: /sn:0 {0}(243,200)(178,200)(178,60)(100,60)(100,19){1}
wire [31:0] R3;    //: {0}(687,228)(687,416){1}
wire [31:0] R1;    //: {0}(281,223)(281,308)(53,308)(53,353){1}
wire w2;    //: /sn:0 {0}(243,212)(204,212){1}
wire [1:0] w11;    //: /sn:0 {0}(-27,-33)(-27,-23)(106,-23)(106,-10){1}
wire [31:0] R0;    //: {0}(77,228)(77,299)(41,299)(41,353){1}
wire [31:0] w5;    //: /sn:0 {0}(675,416)(675,372)(497,372)(497,228){1}
wire [31:0] w9;    //: /sn:0 {0}(663,416)(663,387)(309,387)(309,223){1}
//: enddecls

  //: joint g44 (clr) @(353, -83) /w:[ 3 -1 4 10 ]
  //: input g4 (Read2) @(-239,145) /sn:0 /w:[ 0 ]
  //: joint g8 (w18) @(6, 122) /w:[ 7 -1 8 10 ]
  //: joint g47 (clr) @(541, -83) /w:[ 1 -1 2 12 ]
  //: joint g16 (clk) @(165, 285) /w:[ 5 6 8 -1 ]
  //: input g3 (Write) @(-240,-38) /sn:0 /w:[ 0 ]
  //: joint g26 (w19) @(229, 106) /w:[ 5 -1 6 12 ]
  //: input g17 (Read1) @(-239,96) /sn:0 /w:[ 0 ]
  //: output g2 (Data2) @(668,482) /sn:0 /R:3 /w:[ 0 ]
  tran g30(.Z(w10), .I(Read2[4:3]));   //: @(-140,143) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  tran g23(.Z(w24), .I(Write[2:0]));   //: @(-65,-39) /sn:0 /R:1 /w:[ 9 1 2 ] /ss:1
  Regs8x32 g24 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w31), .clk(w2), .clr(clr), .AOUT(R1), .BOUT(w9));   //: @(244, 153) /sz:(98, 69) /sn:0 /p:[ Ti0>11 Li0>13 Li1>13 Li2>13 Li3>0 Li4>0 Ri0>11 Bo0<0 Bo1<1 ]
  //: joint g39 (RegWrite) @(372, 263) /w:[ 6 8 5 -1 ]
  //: output g1 (Data1) @(59,462) /sn:0 /R:3 /w:[ 1 ]
  Regs8x32 g29 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w4), .clk(w22), .clr(clr), .AOUT(R2), .BOUT(w5));   //: @(432, 158) /sz:(98, 69) /sn:0 /p:[ Ti0>13 Li0>0 Li1>0 Li2>0 Li3>1 Li4>1 Ri0>13 Bo0<1 Bo1<1 ]
  //: comment g51 /dolink:0 /link:"" @(395,229) /sn:0
  //: /line:"Regs 16-23"
  //: /end
  tran g18(.Z(w19), .I(Read1[2:0]));   //: @(-95,93) /sn:0 /R:1 /w:[ 9 3 4 ] /ss:1
  //: joint g25 (w18) @(210, 122) /w:[ 5 -1 6 12 ]
  //: supply1 g10 (w21) @(68,-11) /sn:0 /w:[ 1 ]
  //: comment g49 /dolink:0 /link:"" @(210,225) /sn:0
  //: /line:"Regs 8-15"
  //: /end
  Regs8x32 g6 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w16), .clk(w1), .clr(clr), .AOUT(R0), .BOUT(w0));   //: @(40, 158) /sz:(98, 69) /sn:0 /p:[ Ti0>9 Li0>11 Li1>11 Li2>11 Li3>0 Li4>1 Ri0>9 Bo0<0 Bo1<1 ]
  //: comment g50 /dolink:0 /link:"" @(585,229) /sn:0
  //: /line:"Regs 24-31"
  //: /end
  and g35 (.I0(clk), .I1(RegWrite), .Z(w22));   //: @(394,217) /sn:0 /delay:" 1" /w:[ 3 9 0 ]
  demux g9 (.I(w11), .E(w21), .Z0(w16), .Z1(w31), .Z2(w4), .Z3(w20));   //: @(106,3) /sn:0 /w:[ 1 0 1 1 0 0 ]
  //: joint g7 (w19) @(23, 106) /w:[ 7 -1 8 10 ]
  tran g22(.Z(w18), .I(Read2[2:0]));   //: @(-93,142) /sn:0 /R:1 /w:[ 9 3 4 ] /ss:0
  tran g31(.Z(w6), .I(Read1[4:3]));   //: @(-123,93) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  and g33 (.I0(clk), .I1(RegWrite), .Z(w1));   //: @(-27,217) /sn:0 /delay:" 1" /w:[ 11 13 0 ]
  //: joint g45 (WriteData) @(479, 75) /w:[ 1 -1 2 12 ]
  //: joint g41 (w19) @(419, 107) /w:[ 2 -1 4 1 ]
  and g36 (.I0(clk), .I1(RegWrite), .Z(w23));   //: @(567,217) /sn:0 /delay:" 1" /w:[ 0 7 0 ]
  //: joint g40 (w18) @(402, 123) /w:[ 2 -1 4 1 ]
  //: input g42 (clr) @(-237,-92) /sn:0 /w:[ 7 ]
  //: input g12 (clk) @(-239,285) /sn:0 /w:[ 13 ]
  Regs8x32 g46 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w20), .clk(w23), .clr(clr), .AOUT(w3), .BOUT(R3));   //: @(622, 158) /sz:(98, 69) /sn:0 /p:[ Ti0>0 Li0>3 Li1>3 Li2>3 Li3>1 Li4>1 Ri0>0 Bo0<1 Bo1<0 ]
  //: joint g28 (w24) @(381, 139) /w:[ 2 -1 4 1 ]
  and g34 (.I0(clk), .I1(RegWrite), .Z(w2));   //: @(194,212) /sn:0 /delay:" 1" /w:[ 7 11 1 ]
  tran g5(.Z(w11), .I(Write[4:3]));   //: @(-27,-39) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  mux g14 (.I0(R0), .I1(R1), .I2(R2), .I3(w3), .S(w6), .Z(Data1));   //: @(59,369) /sn:0 /w:[ 1 1 0 0 0 0 ] /ss:0 /do:0
  //: joint g11 (w24) @(-15, 138) /w:[ 7 -1 8 10 ]
  //: joint g21 (w24) @(193, 138) /w:[ 5 -1 6 12 ]
  //: joint g19 (clk) @(-58, 285) /w:[ 9 10 12 -1 ]
  //: joint g20 (WriteData) @(87, 75) /w:[ 5 -1 6 8 ]
  //: input g32 (RegWrite) @(-239,263) /sn:0 /w:[ 0 ]
  //: input g0 (WriteData) @(-239,73) /sn:0 /w:[ 7 ]
  //: joint g43 (clr) @(148, -83) /w:[ 5 -1 6 8 ]
  //: joint g15 (clk) @(362, 285) /w:[ 1 2 4 -1 ]
  //: joint g38 (RegWrite) @(173, 263) /w:[ 4 10 3 -1 ]
  //: comment g48 /dolink:0 /link:"" @(11,228) /sn:0
  //: /line:"Regs 0-7"
  //: /end
  //: joint g27 (WriteData) @(290, 75) /w:[ 3 -1 4 10 ]
  //: joint g37 (RegWrite) @(-69, 263) /w:[ 2 12 1 -1 ]
  mux g13 (.I0(w0), .I1(w9), .I2(w5), .I3(R3), .S(w10), .Z(Data2));   //: @(669,432) /sn:0 /w:[ 0 0 0 1 1 1 ] /ss:0 /do:0

endmodule

module Regs8x32(SB, SA, BOUT, AOUT, clr, clk, RegWr, SD, DIN);
//: interface  /sz:(98, 69) /bd:[ Ti0>DIN[31:0](47/98) Ti1>DIN[31:0](47/98) Ti2>DIN[31:0](47/98) Ti3>DIN[31:0](47/98) Ti4>DIN[31:0](47/98) Ti5>DIN[31:0](47/98) Ti6>DIN[31:0](47/98) Ti7>DIN[31:0](47/98) Ti8>DIN[31:0](47/98) Li0>SD[2:0](35/69) Li1>SA[2:0](11/69) Li2>SB[2:0](22/69) Li3>RegWr(47/69) Li4>clk(59/69) Li5>clk(59/69) Li6>RegWr(47/69) Li7>SB[2:0](22/69) Li8>SA[2:0](11/69) Li9>SD[2:0](35/69) Li10>SD[2:0](35/69) Li11>SA[2:0](11/69) Li12>SB[2:0](22/69) Li13>RegWr(47/69) Li14>clk(59/69) Li15>SD[2:0](35/69) Li16>SA[2:0](11/69) Li17>SB[2:0](22/69) Li18>RegWr(47/69) Li19>clk(59/69) Li20>clk(59/69) Li21>RegWr(47/69) Li22>SB[2:0](22/69) Li23>SA[2:0](11/69) Li24>SD[2:0](35/69) Li25>SD[2:0](35/69) Li26>SA[2:0](11/69) Li27>SB[2:0](22/69) Li28>RegWr(47/69) Li29>clk(59/69) Li30>SD[2:0](35/69) Li31>SA[2:0](11/69) Li32>SB[2:0](22/69) Li33>RegWr(47/69) Li34>clk(59/69) Li35>clk(59/69) Li36>RegWr(47/69) Li37>SB[2:0](22/69) Li38>SA[2:0](11/69) Li39>SD[2:0](35/69) Li40>SD[2:0](35/69) Li41>SA[2:0](11/69) Li42>SB[2:0](22/69) Li43>RegWr(47/69) Li44>clk(59/69) Ri0>clr(35/69) Ri1>clr(35/69) Ri2>clr(35/69) Ri3>clr(35/69) Ri4>clr(35/69) Ri5>clr(35/69) Ri6>clr(35/69) Ri7>clr(35/69) Ri8>clr(35/69) Bo0<AOUT[31:0](37/98) Bo1<BOUT[31:0](65/98) Bo2<BOUT[31:0](65/98) Bo3<AOUT[31:0](37/98) Bo4<AOUT[31:0](37/98) Bo5<BOUT[31:0](65/98) Bo6<AOUT[31:0](37/98) Bo7<BOUT[31:0](65/98) Bo8<BOUT[31:0](65/98) Bo9<AOUT[31:0](37/98) Bo10<AOUT[31:0](37/98) Bo11<BOUT[31:0](65/98) Bo12<AOUT[31:0](37/98) Bo13<BOUT[31:0](65/98) Bo14<BOUT[31:0](65/98) Bo15<AOUT[31:0](37/98) Bo16<AOUT[31:0](37/98) Bo17<BOUT[31:0](65/98) ]
input [31:0] DIN;    //: /sn:0 {0}(531,269)(531,318){1}
//: {2}(533,320)(627,320){3}
//: {4}(631,320)(715,320){5}
//: {6}(719,320)(807,320)(807,429){7}
//: {8}(717,322)(717,352){9}
//: {10}(629,322)(629,433){11}
//: {12}(529,320)(435,320){13}
//: {14}(431,320)(342,320){15}
//: {16}(338,320)(264,320){17}
//: {18}(260,320)(181,320)(181,352){19}
//: {20}(262,322)(262,439){21}
//: {22}(340,322)(340,351){23}
//: {24}(433,322)(433,436){25}
//: {26}(531,322)(531,348){27}
output [31:0] BOUT;    //: /sn:0 {0}(516,697)(516,672){1}
input [2:0] SD;    //: /sn:0 {0}(782,138)(852,138)(852,156){1}
input [2:0] SB;    //: /sn:0 {0}(466,659)(493,659){1}
supply1 w21;    //: /sn:0 {0}(828,169)(801,169)(801,153){1}
input RegWr;    //: /sn:0 {0}(48,363)(68,363)(68,378)(82,378){1}
input clr;    //: /sn:0 /dp:1 {0}(959,337)(1032,337){1}
input [2:0] SA;    //: /sn:0 {0}(256,657)(231,657){1}
input clk;    //: /sn:0 {0}(82,383)(68,383)(68,398)(55,398){1}
output [31:0] AOUT;    //: /sn:0 {0}(279,670)(279,702){1}
wire [31:0] w16;    //: /sn:0 {0}(531,369)(531,574)(520,574){1}
//: {2}(516,574)(282,574)(282,641){3}
//: {4}(518,576)(518,587)(519,587)(519,643){5}
wire w7;    //: /sn:0 {0}(472,451)(513,451)(513,405)(848,405)(848,185){1}
wire [31:0] R5;    //: {0}(288,641)(288,586)(525,586){1}
//: {2}(529,586)(629,586)(629,454){3}
//: {4}(527,588)(527,617)(525,617)(525,643){5}
wire w4;    //: /sn:0 {0}(943,337)(906,337){1}
//: {2}(902,337)(767,337){3}
//: {4}(763,337)(588,337){5}
//: {6}(584,337)(390,337){7}
//: {8}(386,337)(231,337)(231,357)(220,357){9}
//: {10}(388,339)(388,356)(379,356){11}
//: {12}(586,339)(586,353)(570,353){13}
//: {14}(765,339)(765,357)(756,357){15}
//: {16}(904,339)(904,417)(865,417){17}
//: {18}(861,417)(675,417){19}
//: {20}(671,417)(489,417){21}
//: {22}(485,417)(302,417)(302,444)(301,444){23}
//: {24}(487,419)(487,441)(472,441){25}
//: {26}(673,419)(673,438)(668,438){27}
//: {28}(863,419)(863,434)(846,434){29}
wire w3;    //: /sn:0 {0}(835,185)(835,397)(330,397)(330,454)(301,454){1}
wire w0;    //: /sn:0 {0}(770,439)(764,439)(764,481)(579,481){1}
//: {2}(577,479)(577,443)(592,443){3}
//: {4}(575,481)(390,481){5}
//: {6}(388,479)(388,446)(396,446){7}
//: {8}(386,481)(214,481){9}
//: {10}(212,479)(212,449)(225,449){11}
//: {12}(210,481)(125,481)(125,383){13}
//: {14}(127,381)(291,381){15}
//: {16}(295,381)(477,381){17}
//: {18}(481,381)(660,381)(660,362)(680,362){19}
//: {20}(479,379)(479,358)(494,358){21}
//: {22}(293,379)(293,361)(303,361){23}
//: {24}(125,379)(125,362)(144,362){25}
//: {26}(123,381)(103,381){27}
wire [31:0] R2;    //: {0}(262,641)(262,537){1}
//: {2}(264,535)(499,535)(499,643){3}
//: {4}(262,533)(262,460){5}
wire [31:0] R7;    //: {0}(807,450)(807,609)(541,609){1}
//: {2}(537,609)(302,609)(302,641){3}
//: {4}(539,611)(539,643){5}
wire w12;    //: /sn:0 {0}(756,367)(787,367)(787,258)(868,258)(868,185){1}
wire w10;    //: /sn:0 {0}(846,444)(875,444)(875,185){1}
wire [31:0] R4;    //: {0}(340,372)(340,545){1}
//: {2}(342,547)(505,547)(505,643){3}
//: {4}(338,547)(268,547)(268,641){5}
wire [31:0] R3;    //: {0}(512,643)(512,559)(435,559){1}
//: {2}(433,557)(433,457){3}
//: {4}(431,559)(275,559)(275,641){5}
wire w8;    //: /sn:0 {0}(220,367)(249,367)(249,213)(828,213)(828,185){1}
wire Z5;    //: /sn:0 {0}(861,185)(861,413)(700,413)(700,448)(668,448){1}
wire w14;    //: /sn:0 {0}(379,366)(414,366)(414,229)(841,229)(841,185){1}
wire [31:0] R0;    //: {0}(492,643)(492,523)(257,523){1}
//: {2}(253,523)(181,523)(181,373){3}
//: {4}(255,525)(255,641){5}
wire w15;    //: /sn:0 {0}(570,363)(608,363)(608,244)(855,244)(855,185){1}
wire [31:0] R10;    //: /sn:0 {0}(295,641)(295,600)(530,600){1}
//: {2}(534,600)(717,600)(717,373){3}
//: {4}(532,602)(532,643){5}
//: enddecls

  //: input g4 (SB) @(464,659) /sn:0 /w:[ 0 ]
  //: joint g8 (w16) @(518, 574) /w:[ 1 -1 2 4 ]
  //: joint g16 (R3) @(433, 559) /w:[ 1 2 4 -1 ]
  //: input g3 (SA) @(229,657) /sn:0 /w:[ 1 ]
  //: joint g26 (DIN) @(340, 320) /w:[ 15 -1 16 22 ]
  //: joint g17 (R4) @(340, 547) /w:[ 2 1 4 -1 ]
  //: output g2 (BOUT) @(516,694) /sn:0 /R:3 /w:[ 0 ]
  register R5 (.Q(R5), .D(DIN), .EN(Z5), .CLR(w4), .CK(!w0));   //: @(629,443) /w:[ 3 11 1 27 3 ]
  //: joint g30 (w0) @(212, 481) /w:[ 9 10 12 -1 ]
  //: joint g23 (w4) @(765, 337) /w:[ 3 -1 4 14 ]
  //: joint g24 (DIN) @(531, 320) /w:[ 2 1 12 26 ]
  //: joint g39 (DIN) @(262, 320) /w:[ 17 -1 18 20 ]
  //: output g1 (AOUT) @(279,699) /sn:0 /R:3 /w:[ 1 ]
  //: joint g29 (w0) @(388, 481) /w:[ 5 6 8 -1 ]
  register R2 (.Q(R4), .D(DIN), .EN(w14), .CLR(w4), .CK(!w0));   //: @(340,361) /w:[ 0 23 0 11 23 ]
  //: joint g18 (R2) @(262, 535) /w:[ 2 4 -1 1 ]
  register R7 (.Q(R7), .D(DIN), .EN(w10), .CLR(w4), .CK(!w0));   //: @(807,439) /w:[ 0 7 0 29 0 ]
  not g25 (.I(clr), .Z(w4));   //: @(953,337) /sn:0 /R:2 /w:[ 0 0 ]
  //: supply1 g10 (w21) @(812,153) /sn:0 /w:[ 1 ]
  register R6 (.Q(R10), .D(DIN), .EN(w12), .CLR(w4), .CK(!w0));   //: @(717,362) /w:[ 3 9 0 15 19 ]
  //: joint g6 (R7) @(539, 609) /w:[ 1 -1 2 4 ]
  and g35 (.I0(RegWr), .I1(clk), .Z(w0));   //: @(93,381) /sn:0 /delay:" 1" /w:[ 1 0 27 ]
  demux g9 (.I(SD), .E(w21), .Z0(!w8), .Z1(!w3), .Z2(!w14), .Z3(!w7), .Z4(!w15), .Z5(!Z5), .Z6(!w12), .Z7(!w10));   //: @(852,169) /sn:0 /w:[ 1 0 1 0 1 1 1 0 1 1 ]
  register R4 (.Q(w16), .D(DIN), .EN(w15), .CLR(w4), .CK(!w0));   //: @(531,358) /w:[ 0 27 0 13 21 ]
  //: joint g7 (R10) @(532, 600) /w:[ 2 -1 1 4 ]
  //: joint g22 (w4) @(586, 337) /w:[ 5 -1 6 12 ]
  //: joint g31 (w4) @(863, 417) /w:[ 17 -1 18 28 ]
  register R1 (.Q(R2), .D(DIN), .EN(w3), .CLR(w4), .CK(!w0));   //: @(262,449) /w:[ 5 21 1 23 11 ]
  register R3 (.Q(R3), .D(DIN), .EN(w7), .CLR(w4), .CK(!w0));   //: @(433,446) /w:[ 3 25 0 25 7 ]
  //: joint g33 (w4) @(673, 417) /w:[ 19 -1 20 26 ]
  //: joint g41 (DIN) @(717, 320) /w:[ 6 -1 5 8 ]
  //: joint g36 (w4) @(904, 337) /w:[ 1 -1 2 16 ]
  //: joint g40 (DIN) @(433, 320) /w:[ 13 -1 14 24 ]
  //: joint g42 (DIN) @(629, 320) /w:[ 4 -1 3 10 ]
  //: joint g12 (w0) @(479, 381) /w:[ 18 20 17 -1 ]
  //: input g28 (clr) @(1034,337) /sn:0 /R:2 /w:[ 1 ]
  //: input g34 (clk) @(53,398) /sn:0 /w:[ 1 ]
  mux g14 (.I0(R0), .I1(R2), .I2(R4), .I3(R3), .I4(w16), .I5(R5), .I6(R10), .I7(R7), .S(SA), .Z(AOUT));   //: @(279,657) /sn:0 /w:[ 5 0 5 5 3 0 0 3 0 0 ] /ss:0 /do:0
  //: input g5 (RegWr) @(46,363) /sn:0 /w:[ 0 ]
  //: joint g11 (w0) @(293, 381) /w:[ 16 22 15 -1 ]
  //: joint g21 (w4) @(388, 337) /w:[ 7 -1 8 10 ]
  //: joint g19 (R0) @(255, 523) /w:[ 1 -1 2 4 ]
  //: input g20 (SD) @(780,138) /sn:0 /w:[ 0 ]
  //: joint g32 (w4) @(487, 417) /w:[ 21 -1 22 24 ]
  register R0 (.Q(R0), .D(DIN), .EN(w8), .CLR(w4), .CK(!w0));   //: @(181,362) /w:[ 3 19 0 9 25 ]
  //: input g0 (DIN) @(531,267) /sn:0 /R:3 /w:[ 0 ]
  //: joint g15 (R5) @(527, 586) /w:[ 2 -1 1 4 ]
  //: joint g38 (w0) @(577, 481) /w:[ 1 2 4 -1 ]
  //: joint g27 (w0) @(125, 381) /w:[ 14 24 26 13 ]
  mux g13 (.I0(R0), .I1(R2), .I2(R4), .I3(R3), .I4(w16), .I5(R5), .I6(R10), .I7(R7), .S(SB), .Z(BOUT));   //: @(516,659) /sn:0 /w:[ 0 3 3 0 5 5 5 5 1 1 ] /ss:0 /do:0

endmodule

module Read(clk, Inm32, Inst, rs, RegDst, WriteData, clr, rt, RegWrite);
//: interface  /sz:(166, 219) /bd:[ Ti0>RegWrite(84/166) Li0>Inst[31:0](30/219) Li1>RegDst(121/219) Bi0>WriteData[31:0](40/166) Bi1>clr(123/166) Bi2>clk(93/166) Ro0<rs[31:0](51/219) Ro1<rt[31:0](92/219) Ro2<Inm32[31:0](141/219) ]
output [31:0] Inm32;    //: /sn:0 /dp:1 {0}(484,464)(614,464){1}
input [31:0] WriteData;    //: /sn:0 /dp:1 {0}(389,297)(365,297)(365,319)(145,319){1}
output [31:0] rt;    //: /sn:0 /dp:1 {0}(538,288)(627,288){1}
input [31:0] Inst;    //: /sn:0 {0}(212,308)(212,298){1}
//: {2}(212,297)(212,268){3}
//: {4}(212,267)(212,221){5}
//: {6}(212,220)(212,181){7}
//: {8}(212,180)(212,138){9}
input RegDst;    //: /sn:0 {0}(146,348)(318,348)(318,281){1}
input clr;    //: /sn:0 {0}(406,77)(462,77)(462,148){1}
input RegWrite;    //: /sn:0 {0}(145,375)(430,375)(430,332){1}
input clk;    //: /sn:0 {0}(144,397)(498,397)(498,376){1}
output [31:0] rs;    //: /sn:0 {0}(622,196)(538,196){1}
wire [4:0] w6;    //: /sn:0 {0}(216,268)(302,268){1}
wire [4:0] w3;    //: /sn:0 {0}(216,181)(389,181){1}
wire [4:0] w0;    //: /sn:0 {0}(302,248)(262,248)(262,223){1}
//: {2}(264,221)(389,221){3}
//: {4}(260,221)(216,221){5}
wire [4:0] w10;    //: /sn:0 {0}(331,258)(389,258){1}
wire [15:0] w8;    //: /sn:0 /dp:1 {0}(442,462)(224,462)(224,298)(216,298){1}
wire w2;    //: /sn:0 {0}(498,360)(498,332){1}
//: enddecls

  //: joint g4 (w0) @(262, 221) /w:[ 2 -1 4 1 ]
  //: input g8 (clk) @(142,397) /sn:0 /w:[ 0 ]
  mux g3 (.I0(w0), .I1(w6), .S(RegDst), .Z(w10));   //: @(318,258) /sn:0 /R:1 /w:[ 0 1 1 0 ] /ss:0 /do:1
  //: output g16 (Inm32) @(611,464) /sn:0 /w:[ 1 ]
  //: input g17 (Inst) @(212,136) /sn:0 /R:3 /w:[ 9 ]
  tran g2(.Z(w0), .I(Inst[20:16]));   //: @(210,221) /sn:0 /R:2 /w:[ 5 5 6 ] /ss:1
  tran g1(.Z(w3), .I(Inst[25:21]));   //: @(210,181) /sn:0 /R:2 /w:[ 0 7 8 ] /ss:1
  //: output g10 (rs) @(619,196) /sn:0 /w:[ 0 ]
  //: input g6 (RegDst) @(144,348) /sn:0 /w:[ 0 ]
  //: input g7 (WriteData) @(143,319) /sn:0 /w:[ 1 ]
  //: input g9 (clr) @(404,77) /sn:0 /w:[ 0 ]
  not g12 (.I(clk), .Z(w2));   //: @(498,370) /sn:0 /R:1 /w:[ 1 0 ]
  tran g14(.Z(w8), .I(Inst[15:0]));   //: @(210,298) /sn:0 /R:2 /w:[ 1 1 2 ] /ss:1
  tran g5(.Z(w6), .I(Inst[15:11]));   //: @(210,268) /sn:0 /R:2 /w:[ 0 3 4 ] /ss:1
  //: output g11 (rt) @(624,288) /sn:0 /w:[ 1 ]
  BRegs32x32 g0 (.clr(clr), .Read1(w3), .Read2(w0), .Write(w10), .WriteData(WriteData), .clk(w2), .RegWrite(RegWrite), .Data1(rs), .Data2(rt));   //: @(390, 149) /sz:(147, 182) /sn:0 /p:[ Ti0>1 Li0>1 Li1>3 Li2>1 Li3>0 Bi0>1 Bi1>1 Ro0<1 Ro1<0 ]
  Extend g15 (.A(w8), .S(Inm32));   //: @(443, 447) /sz:(40, 40) /sn:0 /p:[ Li0>0 Ro0<0 ]
  //: input g13 (RegWrite) @(143,375) /sn:0 /w:[ 0 ]

endmodule

module Extend(S, A);
//: interface  /sz:(40, 40) /bd:[ Li0>A[15:0](23/40) Li1>A[15:0](23/40) Ro0<S[31:0](23/40) Ro1<S[31:0](23/40) ]
input [15:0] A;    //: /sn:0 {0}(307,243)(307,412)(325,412){1}
//: {2}(326,412)(355,412){3}
output [31:0] S;    //: /sn:0 /dp:1 {0}(361,332)(401,332){1}
wire w1;    //: /sn:0 {0}(326,407)(326,404){1}
//: {2}(328,402)(355,402){3}
//: {4}(326,400)(326,394){5}
//: {6}(328,392)(355,392){7}
//: {8}(326,390)(326,384){9}
//: {10}(328,382)(355,382){11}
//: {12}(326,380)(326,374){13}
//: {14}(328,372)(355,372){15}
//: {16}(326,370)(326,364){17}
//: {18}(328,362)(355,362){19}
//: {20}(326,360)(326,354){21}
//: {22}(328,352)(355,352){23}
//: {24}(326,350)(326,344){25}
//: {26}(328,342)(355,342){27}
//: {28}(326,340)(326,334){29}
//: {30}(328,332)(355,332){31}
//: {32}(326,330)(326,324){33}
//: {34}(328,322)(355,322){35}
//: {36}(326,320)(326,314){37}
//: {38}(328,312)(355,312){39}
//: {40}(326,310)(326,304){41}
//: {42}(328,302)(355,302){43}
//: {44}(326,300)(326,294){45}
//: {46}(328,292)(355,292){47}
//: {48}(326,290)(326,284){49}
//: {50}(328,282)(355,282){51}
//: {52}(326,280)(326,274){53}
//: {54}(328,272)(355,272){55}
//: {56}(326,270)(326,264){57}
//: {58}(328,262)(355,262){59}
//: {60}(326,260)(326,252)(355,252){61}
//: enddecls

  //: joint g8 (w1) @(326, 382) /w:[ 10 12 -1 9 ]
  tran g4(.Z(w1), .I(A[15]));   //: @(326,410) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:0
  //: joint g16 (w1) @(326, 302) /w:[ 42 44 -1 41 ]
  //: joint g17 (w1) @(326, 292) /w:[ 46 48 -1 45 ]
  concat g2 (.I0(A), .I1(w1), .I2(w1), .I3(w1), .I4(w1), .I5(w1), .I6(w1), .I7(w1), .I8(w1), .I9(w1), .I10(w1), .I11(w1), .I12(w1), .I13(w1), .I14(w1), .I15(w1), .I16(w1), .Z(S));   //: @(360,332) /sn:0 /w:[ 3 3 7 11 15 19 23 27 31 35 39 43 47 51 55 59 61 0 ] /dr:0
  //: output g1 (S) @(398,332) /sn:0 /w:[ 1 ]
  //: joint g18 (w1) @(326, 282) /w:[ 50 52 -1 49 ]
  //: joint g10 (w1) @(326, 362) /w:[ 18 20 -1 17 ]
  //: joint g9 (w1) @(326, 372) /w:[ 14 16 -1 13 ]
  //: joint g7 (w1) @(326, 392) /w:[ 6 8 -1 5 ]
  //: joint g12 (w1) @(326, 342) /w:[ 26 28 -1 25 ]
  //: joint g14 (w1) @(326, 322) /w:[ 34 36 -1 33 ]
  //: joint g11 (w1) @(326, 352) /w:[ 22 24 -1 21 ]
  //: joint g5 (w1) @(326, 402) /w:[ 2 4 -1 1 ]
  //: joint g19 (w1) @(326, 272) /w:[ 54 56 -1 53 ]
  //: joint g20 (w1) @(326, 262) /w:[ 58 60 -1 57 ]
  //: joint g15 (w1) @(326, 312) /w:[ 38 40 -1 37 ]
  //: input g0 (A) @(307,241) /sn:0 /R:3 /w:[ 0 ]
  //: joint g13 (w1) @(326, 332) /w:[ 30 32 -1 29 ]

endmodule

module main;    //: root_module
wire w13;    //: /sn:0 {0}(1365,410)(1365,137)(778,137){1}
wire [31:0] w6;    //: /sn:0 /dp:5 {0}(834,442)(724,442)(724,482){1}
//: {2}(724,483)(724,513){3}
//: {4}(724,514)(724,564)(680,564){5}
wire [31:0] w16;    //: /sn:0 /dp:1 {0}(1163,303)(1279,303)(1279,321)(1315,321){1}
wire [31:0] w7;    //: /sn:0 {0}(680,449)(692,449)(692,331)(1010,331){1}
//: {2}(1014,331)(1028,331){3}
//: {4}(1029,331)(1234,331){5}
//: {6}(1012,333)(1012,438)(1041,438){7}
wire Zero;    //: /sn:0 /dp:1 {0}(1185,444)(1213,444)(1213,246)(1248,246)(1248,256){1}
wire w4;    //: /sn:0 {0}(590,571)(523,571)(523,863){1}
//: {2}(525,865)(909,865){3}
//: {4}(913,865)(1500,865){5}
//: {6}(911,863)(911,632){7}
//: {8}(521,865)(483,865){9}
wire [31:0] Inm32;    //: /sn:0 /dp:1 {0}(973,561)(1041,561){1}
wire w0;    //: /sn:0 {0}(1465,484)(1465,118)(778,118){1}
wire [31:0] w3;    //: /sn:0 /dp:3 {0}(1478,507)(1526,507)(1526,693)(868,693)(868,665){1}
//: {2}(868,664)(868,632){3}
wire w20;    //: /sn:0 {0}(778,69)(1331,69)(1331,308){1}
wire [31:0] rt;    //: /sn:0 /dp:1 {0}(1041,527)(1018,527){1}
//: {2}(1014,527)(973,527){3}
//: {4}(1016,529)(1016,633)(1196,633)(1196,559)(1253,559){5}
wire w19;    //: /sn:0 {0}(778,84)(1253,84)(1253,256){1}
wire [31:0] w12;    //: /sn:0 {0}(1185,462)(1199,462)(1199,351)(1234,351){1}
wire [3:0] w23;    //: /sn:0 /dp:1 {0}(778,226)(1093,226)(1093,377)(1129,377)(1129,412){1}
wire w10;    //: /sn:0 /dp:1 {0}(1250,318)(1250,277){1}
wire [31:0] ALUResult;    //: /sn:0 /dp:1 {0}(1185,488)(1227,488){1}
//: {2}(1231,488)(1253,488){3}
//: {4}(1229,490)(1229,644)(1432,644)(1432,517)(1449,517){5}
wire w21;    //: /sn:0 {0}(1294,410)(1294,102)(778,102){1}
wire [31:0] w1;    //: /sn:0 {0}(1449,497)(1425,497)(1425,489)(1402,489){1}
wire RegDst;    //: /sn:0 {0}(834,533)(788,533)(788,261)(778,261){1}
wire [25:0] w8;    //: /sn:0 {0}(863,665)(753,665)(753,308)(1157,308){1}
wire w27;    //: /sn:0 {0}(778,172)(904,172)(904,411){1}
wire [5:0] w17;    //: /sn:0 {0}(728,514)(737,514)(737,284){1}
wire [31:0] w14;    //: /sn:0 /dp:1 {0}(1344,331)(1503,331)(1503,40)(582,40)(582,424)(590,424){1}
wire [31:0] w11;    //: /sn:0 /dp:1 {0}(1263,341)(1315,341){1}
wire w2;    //: /sn:0 {0}(936,751)(936,632){1}
wire [5:0] w15;    //: /sn:0 {0}(1029,326)(1029,298)(1157,298){1}
wire [5:0] w5;    //: /sn:0 {0}(719,483)(710,483)(710,284){1}
wire w26;    //: /sn:0 {0}(778,153)(1068,153)(1068,412){1}
wire w9;    //: /sn:0 {0}(522,455)(590,455){1}
wire [31:0] rs;    //: /sn:0 {0}(1041,494)(973,494){1}
//: enddecls

  //: joint g8 (w4) @(523, 865) /w:[ 2 1 8 -1 ]
  mux g4 (.I0(ALUResult), .I1(w1), .S(w0), .Z(w3));   //: @(1465,507) /sn:0 /R:1 /w:[ 5 0 0 0 ] /ss:1 /do:0
  Mem g3 (.MemRead(w21), .MemWrite(w13), .WriteData(rt), .Adress(ALUResult), .ReadData(w1));   //: @(1254, 411) /sz:(147, 210) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>5 Li1>3 Ro0<1 ]
  tran g16(.Z(w15), .I(w7[31:26]));   //: @(1029,329) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:0
  //: comment g17 /dolink:0 /link:"" @(1319,280) /sn:0
  //: /line:"Jump"
  //: /end
  //: joint g2 (rt) @(1016, 527) /w:[ 1 -1 2 4 ]
  tran g23(.Z(w17), .I(w6[5:0]));   //: @(722,514) /sn:0 /R:2 /w:[ 0 4 3 ] /ss:1
  and g24 (.I0(w19), .I1(Zero), .Z(w10));   //: @(1250,267) /sn:0 /R:3 /w:[ 1 1 1 ]
  EXE g1 (.ALUSrc(w26), .ALUOperation(w23), .PCNext(w7), .Inm32(Inm32), .rs(rs), .rt(rt), .BranchTarget(w12), .Zero(Zero), .ALUResult(ALUResult));   //: @(1042, 413) /sz:(142, 213) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>7 Li1>1 Li2>0 Li3>0 Ro0<0 Ro1<0 Ro2<0 ]
  //: switch g18 (w2) @(936,765) /sn:0 /R:1 /w:[ 0 ] /st:0
  //: joint g10 (w7) @(1012, 331) /w:[ 2 -1 1 6 ]
  fetch g6 (.Reset(w9), .Clk(w4), .PCNew(w14), .PCNext(w7), .Inst(w6));   //: @(591, 411) /sz:(88, 222) /sn:0 /p:[ Li0>1 Li1>0 Li2>1 Ro0<0 Ro1<5 ]
  //: joint g9 (w4) @(911, 865) /w:[ 4 6 3 -1 ]
  clock g7 (.Z(w4));   //: @(470,865) /sn:0 /w:[ 9 ] /omega:1000 /phi:0 /duty:50
  tran g22(.Z(w5), .I(w6[26:31]));   //: @(722,483) /sn:0 /R:2 /w:[ 0 2 1 ] /ss:0
  //: comment g12 /dolink:0 /link:"" @(1219,282) /sn:0
  //: /line:"PCSrc"
  //: /end
  //: joint g5 (ALUResult) @(1229, 488) /w:[ 2 -1 1 4 ]
  mux g11 (.I0(w7), .I1(w12), .S(w10), .Z(w11));   //: @(1250,341) /sn:0 /R:1 /w:[ 5 1 0 0 ] /ss:1 /do:1
  concat g14 (.I0(w8), .I1(w15), .Z(w16));   //: @(1162,303) /sn:0 /w:[ 1 1 0 ] /dr:0
  UC g21 (.Funct(w17), .Op(w5), .RegDst(RegDst), .RegWrite(w27), .ALUSrc(w26), .MemWrite(w13), .ALUCtrl(w23), .MemToRed(w0), .MemRead(w21), .Jump(w20), .Branch(w19));   //: @(676, 52) /sz:(101, 231) /sn:0 /p:[ Bi0>1 Bi1>1 Ro0<1 Ro1<0 Ro2<0 Ro3<1 Ro4<0 Ro5<1 Ro6<1 Ro7<0 Ro8<0 ]
  //: switch g19 (w9) @(505,455) /sn:0 /w:[ 0 ] /st:0
  //: comment g20 /dolink:0 /link:"" @(1473,465) /sn:0
  //: /line:"MemtoReg"
  //: /end
  Read g0 (.RegWrite(w27), .RegDst(RegDst), .Inst(w6), .clk(w4), .clr(w2), .WriteData(w3), .Inm32(Inm32), .rt(rt), .rs(rs));   //: @(835, 412) /sz:(137, 219) /sn:0 /p:[ Ti0>1 Li0>0 Li1>0 Bi0>7 Bi1>1 Bi2>3 Ro0<0 Ro1<3 Ro2<1 ]
  tran g15(.Z(w8), .I(w3[25:0]));   //: @(866,665) /sn:0 /R:2 /w:[ 0 1 2 ] /ss:0
  mux g13 (.I0(w11), .I1(w16), .S(w20), .Z(w14));   //: @(1331,331) /sn:0 /R:1 /w:[ 1 1 1 0 ] /ss:1 /do:0

endmodule
