//: version "1.8.7"

module fetch(Clk, PCNew, Reset, PCNext, Inst);
//: interface  /sz:(88, 222) /bd:[ Li0>PCNew[31:0](13/222) Li1>Clk(160/222) Li2>Reset(44/222) Ro0<Inst[31:0](159/222) Ro1<PCNext[31:0](38/222) ]
input Clk;    //: /sn:0 {0}(122,387)(184,387)(184,357){1}
input [31:0] PCNew;    //: /sn:0 {0}(124,319)(173,319){1}
output [31:0] Inst;    //: /sn:0 /dp:1 {0}(330,317)(369,317){1}
output [31:0] PCNext;    //: /sn:0 {0}(416,153)(360,153){1}
input Reset;    //: /sn:0 {0}(124,265)(179,265)(179,281){1}
supply0 [31:0] w11;    //: /sn:0 {0}(331,169)(323,169){1}
//: {2}(322,169)(314,169)(314,178){3}
wire Cout;    //: /sn:0 {0}(345,177)(345,187){1}
wire w2;    //: /sn:0 {0}(189,281)(189,153)(212,153){1}
//: {2}(216,153)(323,153)(323,164){3}
//: {4}(214,151)(214,116)(345,116)(345,129){5}
//: {6}(214,155)(214,358)(313,358)(313,344){7}
wire [31:0] x;    //: /sn:0 /dp:4 {0}(194,319)(243,319){1}
//: {2}(247,319)(295,319){3}
//: {4}(245,317)(245,137)(331,137){5}
//: enddecls

  //: input g8 (Clk) @(120,387) /sn:0 /w:[ 0 ]
  //: supply0 g3 (w11) @(314,184) /sn:0 /w:[ 3 ]
  add g2 (.A(w11), .B(x), .S(PCNext), .CI(!w2), .CO(Cout));   //: @(347,153) /sn:0 /R:1 /w:[ 0 5 1 5 0 ]
  register g1 (.Q(x), .D(PCNew), .EN(w2), .CLR(!Reset), .CK(!Clk));   //: @(184,319) /sn:0 /R:1 /w:[ 0 1 0 1 1 ]
  tran g10(.Z(w2), .I(w11[0]));   //: @(323,167) /sn:0 /R:1 /w:[ 3 2 1 ] /ss:0
  //: input g6 (PCNew) @(122,319) /sn:0 /w:[ 0 ]
  //: input g9 (Reset) @(122,265) /sn:0 /w:[ 0 ]
  //: output g7 (PCNext) @(413,153) /sn:0 /w:[ 0 ]
  //: output g12 (Inst) @(366,317) /sn:0 /w:[ 1 ]
  //: joint g5 (x) @(245, 319) /w:[ 2 4 1 -1 ]
  //: joint g11 (w2) @(214, 153) /w:[ 2 4 1 6 ]
  rom g0 (.A(x), .D(Inst), .OE(w2));   //: @(313,318) /sn:0 /w:[ 3 0 7 ] /mem:"/home/milax/Documents/EC/EC_Prac2_V2/mult.mem"

endmodule

module main;    //: root_module
wire Clk;    //: /sn:0 {0}(154,298)(222,298){1}
wire [31:0] PCNew;    //: /sn:0 {0}(519,92)(519,126)(355,126){1}
//: {2}(353,124)(353,53)(214,53)(214,151)(222,151){3}
//: {4}(353,128)(353,176)(312,176){5}
wire [31:0] Inst;    //: /sn:0 {0}(528,249)(528,297)(312,297){1}
wire w1;    //: /sn:0 {0}(178,182)(222,182){1}
//: enddecls

  clock g4 (.Z(Clk));   //: @(141,298) /sn:0 /w:[ 0 ] /omega:600 /phi:0 /duty:50
  //: joint g1 (PCNew) @(353, 126) /w:[ 1 2 -1 4 ]
  led g6 (.I(Inst));   //: @(528,242) /sn:0 /w:[ 0 ] /type:2
  //: switch g9 (w1) @(161,182) /sn:0 /w:[ 0 ] /st:0
  led g7 (.I(PCNew));   //: @(519,85) /sn:0 /w:[ 0 ] /type:2
  fetch g0 (.PCNew(PCNew), .Clk(Clk), .Reset(w1), .Inst(Inst), .PCNext(PCNew));   //: @(223, 138) /sz:(88, 222) /sn:0 /p:[ Li0>3 Li1>1 Li2>1 Ro0<1 Ro1<5 ]

endmodule
