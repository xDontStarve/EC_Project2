//: version "1.8.7"

module UC(ALUCtrl, Func, MemRead, MemToReg, MemWrite, RegWrite, RegDst, ALUSrc, Op, Branch, Jump);
//: interface  /sz:(101, 231) /bd:[ Bi0>Func[5:0](61/101) Bi1>Op[5:0](34/101) Ro0<RegDst(209/231) Ro1<RegWrite(120/231) Ro2<ALUSrc(101/231) Ro3<MemWrite(85/231) Ro4<ALUCtrl[3:0](174/231) Ro5<MemToReg(66/231) Ro6<MemRead(50/231) Ro7<Jump(17/231) Ro8<Branch(32/231) ]
output Branch;    //: /sn:0 /dp:1 {0}(515,270)(678,270){1}
output [3:0] ALUCtrl;    //: /sn:0 /dp:1 {0}(515,163)(672,163){1}
supply0 [31:0] w29;    //: /sn:0 {0}(50,141)(50,145){1}
//: {2}(50,146)(50,156)(35,156)(35,25){3}
//: {4}(37,23)(332,23){5}
//: {6}(333,23)(354,23){7}
//: {8}(35,21)(35,0)(-133,0){9}
//: {10}(-134,0)(-279,0){11}
output MemWrite;    //: /sn:0 /dp:1 {0}(515,141)(674,141){1}
output ALUSrc;    //: /sn:0 /dp:1 {0}(515,116)(673,116){1}
output RegDst;    //: /sn:0 /dp:1 {0}(515,294)(676,294){1}
supply1 w32;    //: /sn:0 {0}(175,127)(175,134){1}
//: {2}(177,136)(275,136){3}
//: {4}(175,138)(175,176)(275,176){5}
output RegWrite;    //: /sn:0 {0}(673,92)(515,92){1}
input [5:0] Op;    //: /sn:0 {0}(152,-93)(152,-70)(367,-70){1}
//: {2}(368,-70)(416,-70){3}
//: {4}(417,-70)(448,-70){5}
input [5:0] Func;    //: /sn:0 {0}(-54,202)(141,202){1}
//: {2}(142,202)(171,202){3}
//: {4}(172,202)(187,202)(187,208){5}
output MemRead;    //: /sn:0 /dp:1 {0}(515,218)(675,218){1}
output MemToReg;    //: /sn:0 /dp:1 {0}(515,193)(672,193){1}
output Jump;    //: /sn:0 /dp:1 {0}(515,247)(674,247){1}
wire [11:0] w13;    //: /sn:0 /dp:1 {0}(471,85)(511,85)(511,91){1}
//: {2}(511,92)(511,115){3}
//: {4}(511,116)(511,140){5}
//: {6}(511,141)(511,162){7}
//: {8}(511,163)(511,192){9}
//: {10}(511,193)(511,217){11}
//: {12}(511,218)(511,246){13}
//: {14}(511,247)(511,269){15}
//: {16}(511,270)(511,293){17}
//: {18}(511,294)(511,312){19}
wire [11:0] w7;    //: /sn:0 {0}(333,27)(333,69){1}
//: {2}(335,71)(352,71){3}
//: {4}(331,71)(329,71){5}
//: {6}(325,71)(316,71)(316,85)(352,85){7}
//: {8}(327,73)(327,78)(352,78){9}
//: {10}(333,73)(333,111)(352,111){11}
wire w25;    //: /sn:0 {0}(172,206)(172,245)(204,245)(204,276){1}
wire [11:0] w4;    //: /sn:0 {0}(238,41)(238,98)(352,98){1}
wire [2:0] w22;    //: /sn:0 {0}(142,206)(142,286){1}
wire [11:0] w0;    //: /sn:0 {0}(188,69)(188,105)(352,105){1}
wire [2:0] w3;    //: /sn:0 {0}(368,-66)(368,72){1}
wire [3:0] w30;    //: /sn:0 /dp:3 {0}(275,146)(72,146){1}
//: {2}(71,146)(54,146){3}
wire [3:0] w18;    //: /sn:0 /dp:1 {0}(188,309)(155,309){1}
wire [3:0] w19;    //: /sn:0 /dp:1 {0}(126,298)(-17,298)(-17,476)(137,476)(137,469){1}
wire w12;    //: /sn:0 {0}(417,-66)(417,-55)(458,-55)(458,62){1}
wire [3:0] w23;    //: /sn:0 {0}(64,251)(64,269)(169,269)(169,289)(188,289){1}
wire [3:0] w10;    //: /sn:0 /dp:1 {0}(136,401)(136,405)(7,405)(7,318)(126,318){1}
wire [3:0] w21;    //: /sn:0 {0}(-133,4)(-133,285)(-80,285){1}
//: {2}(-76,285)(-70,285){3}
//: {4}(-66,285)(-63,285){5}
//: {6}(-59,285)(126,285){7}
//: {8}(-61,287)(-61,292)(126,292){9}
//: {10}(-68,287)(-68,312)(126,312){11}
//: {12}(-78,287)(-78,325)(126,325){13}
wire [3:0] w8;    //: /sn:0 {0}(136,370)(136,374)(17,374)(17,332)(126,332){1}
wire [1:0] w27;    //: /sn:0 {0}(72,150)(72,166)(275,166){1}
wire [11:0] w28;    //: /sn:0 /dp:1 {0}(281,156)(318,156)(318,118)(352,118){1}
wire [11:0] w14;    //: /sn:0 /dp:1 {0}(413,3)(413,75)(442,75){1}
wire [11:0] w2;    //: /sn:0 /dp:1 {0}(300,15)(300,91)(352,91){1}
wire [3:0] w15;    //: /sn:0 {0}(136,432)(136,442)(-4,442)(-4,305)(126,305){1}
wire [3:0] w26;    //: /sn:0 {0}(217,299)(237,299)(237,156)(275,156){1}
wire [11:0] w9;    //: /sn:0 {0}(381,95)(442,95){1}
//: enddecls

  tran g44(.Z(ALUSrc), .I(w13[1]));   //: @(509,116) /sn:0 /R:2 /w:[ 0 4 3 ] /ss:1
  //: comment g8 /dolink:0 /link:"" @(192,71) /sn:0
  //: /line:"Jump"
  //: /end
  //: dip g4 (w0) @(188,59) /sn:0 /w:[ 0 ] /st:512
  //: output g47 (ALUCtrl) @(669,163) /sn:0 /w:[ 1 ]
  //: dip g3 (w8) @(136,360) /sn:0 /w:[ 0 ] /st:2
  //: comment g16 /dolink:0 /link:"" @(430,-37) /sn:0
  //: /line:"SW"
  //: /end
  mux g26 (.I0(w18), .I1(w23), .S(w25), .Z(w26));   //: @(204,299) /sn:0 /R:1 /w:[ 0 1 1 0 ] /ss:1 /do:0
  mux g17 (.I0(w8), .I1(w21), .I2(w10), .I3(w21), .I4(w15), .I5(w19), .I6(w21), .I7(w21), .S(w22), .Z(w18));   //: @(142,309) /sn:0 /R:1 /w:[ 1 13 1 11 1 0 9 7 1 1 ] /ss:1 /do:0
  mux g2 (.I0(w28), .I1(w7), .I2(w0), .I3(w4), .I4(w2), .I5(w7), .I6(w7), .I7(w7), .S(w3), .Z(w9));   //: @(368,95) /sn:0 /R:1 /w:[ 1 11 1 1 1 7 9 3 1 0 ] /ss:1 /do:0
  //: comment g30 /dolink:0 /link:"" @(105,232) /sn:0
  //: /line:"Slt"
  //: /end
  //: comment g23 /dolink:0 /link:"" @(181,380) /sn:0
  //: /line:"Sub"
  //: /end
  //: comment g39 /dolink:0 /link:"" @(106,108) /sn:0
  //: /line:"RegDst & RegWrite active"
  //: /end
  //: comment g24 /dolink:0 /link:"" @(180,412) /sn:0
  //: /line:"And"
  //: /end
  //: input g1 (Func) @(-56,202) /sn:0 /w:[ 0 ]
  //: joint g60 (w29) @(35, 23) /w:[ 4 8 -1 3 ]
  //: dip g29 (w23) @(64,241) /sn:0 /w:[ 0 ] /st:7
  //: output g51 (MemRead) @(672,218) /sn:0 /w:[ 1 ]
  //: dip g18 (w10) @(136,391) /sn:0 /w:[ 0 ] /st:6
  //: joint g65 (w21) @(-61, 285) /w:[ 6 -1 5 8 ]
  //: comment g25 /dolink:0 /link:"" @(181,453) /sn:0
  //: /line:"Or"
  //: /end
  //: comment g10 /dolink:0 /link:"" @(258,80) /sn:0
  //: /line:"lw"
  //: /end
  tran g64(.Z(w21), .I(w29[3:0]));   //: @(-133,-2) /sn:0 /R:1 /w:[ 0 10 9 ] /ss:1
  //: output g49 (MemToReg) @(669,193) /sn:0 /w:[ 1 ]
  tran g50(.Z(MemToReg), .I(w13[7]));   //: @(509,193) /sn:0 /R:2 /w:[ 0 10 9 ] /ss:1
  //: comment g6 /dolink:0 /link:"" @(335,118) /sn:0
  //: /line:"ALU"
  //: /end
  tran g58(.Z(RegDst), .I(w13[11]));   //: @(509,294) /sn:0 /R:2 /w:[ 0 18 17 ] /ss:1
  tran g56(.Z(Branch), .I(w13[10]));   //: @(509,270) /sn:0 /R:2 /w:[ 0 16 15 ] /ss:1
  tran g35(.Z(w27), .I(w30[1:0]));   //: @(72,144) /sn:0 /R:1 /w:[ 0 2 1 ] /ss:1
  //: dip g9 (w4) @(238,31) /sn:0 /w:[ 0 ] /st:403
  //: comment g7 /dolink:0 /link:"" @(308,59) /sn:0
  //: /line:"BEQ"
  //: /end
  //: comment g59 /dolink:0 /link:"" @(-268,-38) /sn:0
  //: /line:"Universal Trash Provider"
  //: /end
  //: comment g31 /dolink:0 /link:"" @(10,173) /sn:0
  //: /line:"Filter add, sub, and & or"
  //: /end
  //: comment g22 /dolink:0 /link:"" @(180,351) /sn:0
  //: /line:"Add"
  //: /end
  //: joint g67 (w21) @(-78, 285) /w:[ 2 -1 1 12 ]
  tran g54(.Z(Jump), .I(w13[9]));   //: @(509,247) /sn:0 /R:2 /w:[ 0 14 13 ] /ss:1
  //: output g45 (MemWrite) @(671,141) /sn:0 /w:[ 1 ]
  //: output g41 (RegWrite) @(670,92) /sn:0 /w:[ 0 ]
  //: supply1 g36 (w32) @(186,127) /sn:0 /w:[ 0 ]
  //: supply0 g33 (w29) @(-285,0) /sn:0 /R:3 /w:[ 11 ]
  tran g52(.Z(MemRead), .I(w13[8]));   //: @(509,218) /sn:0 /R:2 /w:[ 0 12 11 ] /ss:1
  tran g42(.Z(RegWrite), .I(w13[0]));   //: @(509,92) /sn:0 /R:2 /w:[ 1 2 1 ] /ss:1
  //: comment g40 /dolink:0 /link:"" @(113,-43) /sn:0
  //: /line:"OP:"
  //: /line:"   lw: 0010 0011"
  //: /line:"   sw: 0010 1011"
  //: /line:"   beq:0000 0100"
  //: /line:"   j:  0000 0010"
  //: /end
  //: joint g66 (w21) @(-68, 285) /w:[ 4 -1 3 10 ]
  mux g12 (.I0(w9), .I1(w14), .S(w12), .Z(w13));   //: @(458,85) /sn:0 /R:1 /w:[ 1 1 1 0 ] /ss:1 /do:0
  //: output g57 (RegDst) @(673,294) /sn:0 /w:[ 1 ]
  tran g46(.Z(MemWrite), .I(w13[2]));   //: @(509,141) /sn:0 /R:2 /w:[ 0 6 5 ] /ss:1
  tran g34(.Z(w30), .I(w29[3:0]));   //: @(48,146) /sn:0 /R:2 /w:[ 3 2 1 ] /ss:1
  //: comment g28 /dolink:0 /link:"" @(231,310) /sn:0
  //: /line:"Filter whether it's "
  //: /line:"slt or others (bit 3 of func):"
  //: /line:"others: 0010 [0] xxx"
  //: /line:"slt:    0010 [1] 010"
  //: /end
  //: comment g14 /dolink:0 /link:"" @(389,-133) /sn:0
  //: /line:"Determine whether it's SW or others (third bit)"
  //: /line:"LW: 0010 0 011"
  //: /line:"SW: 0010 1 011"
  //: /line:"ALU:0000 0 000"
  //: /end
  tran g11(.Z(w3), .I(Op[2:0]));   //: @(368,-72) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: dip g5 (w2) @(300,5) /sn:0 /w:[ 0 ] /st:1072
  tran g61(.Z(w7), .I(w29[11:0]));   //: @(333,21) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  tran g21(.Z(w22), .I(Func[2:0]));   //: @(142,200) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: dip g19 (w15) @(136,422) /sn:0 /w:[ 0 ] /st:0
  concat g32 (.I0(w32), .I1(w27), .I2(w26), .I3(w30), .I4(w32), .Z(w28));   //: @(280,156) /sn:0 /w:[ 5 1 1 0 3 0 ] /dr:0
  //: dip g20 (w19) @(137,459) /sn:0 /w:[ 1 ] /st:1
  //: joint g63 (w7) @(327, 71) /w:[ 5 -1 6 8 ]
  //: output g43 (ALUSrc) @(670,116) /sn:0 /w:[ 1 ]
  //: comment g38 /dolink:0 /link:"" @(-235,134) /sn:0
  //: /line:"0 value in others signals for ALU instructions"
  //: /end
  //: dip g15 (w14) @(413,-7) /sn:0 /w:[ 0 ] /st:22
  //: input g0 (Op) @(152,-95) /sn:0 /R:3 /w:[ 0 ]
  tran g48(.Z(ALUCtrl), .I(w13[6:3]));   //: @(509,163) /sn:0 /R:2 /w:[ 0 8 7 ] /ss:1
  tran g27(.Z(w25), .I(Func[3]));   //: @(172,200) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  //: joint g62 (w7) @(333, 71) /w:[ 2 1 4 10 ]
  //: joint g37 (w32) @(175, 136) /w:[ 2 1 -1 4 ]
  //: output g55 (Branch) @(675,270) /sn:0 /w:[ 1 ]
  //: output g53 (Jump) @(671,247) /sn:0 /w:[ 1 ]
  tran g13(.Z(w12), .I(Op[3]));   //: @(417,-72) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1

endmodule

module Mem(MemRead, MemWrite, WriteData, ReadData, Address);
//: interface  /sz:(147, 210) /bd:[ Ti0>MemRead(40/147) Ti1>MemWrite(111/147) Li0>WriteData[31:0](148/210) Li1>Address[31:0](77/210) Ro0<ReadData[31:0](78/210) ]
output [31:0] ReadData;    //: /sn:0 /dp:1 {0}(596,161)(660,161){1}
//: {2}(664,161)(854,161){3}
//: {4}(662,163)(662,172){5}
supply0 w0;    //: /sn:0 {0}(572,208)(572,188){1}
input [31:0] WriteData;    //: /sn:0 {0}(740,179)(750,179)(750,194)(662,194)(662,188){1}
input MemWrite;    //: /sn:0 {0}(562,71)(579,71)(579,93){1}
//: {2}(581,95)(636,95)(636,180)(657,180){3}
//: {4}(579,97)(579,138){5}
input MemRead;    //: /sn:0 {0}(529,226)(586,226)(586,188){1}
input [31:0] Address;    //: /sn:0 /dp:1 {0}(561,163)(539,163)(539,130)(334,130){1}
//: enddecls

  //: supply0 g4 (w0) @(572,214) /sn:0 /w:[ 0 ]
  //: joint g8 (ReadData) @(662, 161) /w:[ 2 -1 1 4 ]
  //: input g3 (MemRead) @(527,226) /sn:0 /w:[ 0 ]
  //: input g2 (MemWrite) @(560,71) /sn:0 /w:[ 0 ]
  ram g1 (.A(Address), .D(ReadData), .WE(!MemWrite), .OE(!MemRead), .CS(w0));   //: @(579,162) /sn:0 /w:[ 0 0 5 1 1 ]
  //: joint g10 (MemWrite) @(579, 95) /w:[ 2 1 -1 4 ]
  bufif1 g6 (.Z(ReadData), .I(WriteData), .E(MemWrite));   //: @(662,182) /sn:0 /R:1 /w:[ 5 1 3 ]
  //: input g7 (WriteData) @(738,179) /sn:0 /w:[ 0 ]
  //: output g9 (ReadData) @(851,161) /sn:0 /w:[ 3 ]
  //: comment g5 /dolink:0 /link:"" @(370,188) /sn:0
  //: /line:"Negate to write on low cycle"
  //: /end
  //: input g0 (Address) @(332,130) /sn:0 /w:[ 1 ]

endmodule

module fetch(Clk, PCNew, Reset, PCNext, Inst);
//: interface  /sz:(88, 222) /bd:[ Li0>PCNew[31:0](13/222) Li1>Clk(160/222) Li2>Reset(44/222) Ro0<Inst[31:0](159/222) Ro1<PCNext[31:0](38/222) ]
input Clk;    //: /sn:0 {0}(122,387)(184,387)(184,357){1}
input [31:0] PCNew;    //: /sn:0 {0}(124,319)(173,319){1}
output [31:0] Inst;    //: /sn:0 /dp:1 {0}(330,317)(369,317){1}
output [31:0] PCNext;    //: /sn:0 {0}(416,153)(360,153){1}
input Reset;    //: /sn:0 {0}(124,265)(179,265)(179,281){1}
supply0 [31:0] w11;    //: /sn:0 {0}(331,169)(323,169){1}
//: {2}(322,169)(314,169)(314,178){3}
wire Cout;    //: /sn:0 {0}(345,177)(345,187){1}
wire w2;    //: /sn:0 {0}(189,281)(189,153)(212,153){1}
//: {2}(216,153)(323,153)(323,164){3}
//: {4}(214,151)(214,116)(345,116)(345,129){5}
//: {6}(214,155)(214,358)(313,358)(313,344){7}
wire [31:0] x;    //: /sn:0 /dp:4 {0}(194,319)(243,319){1}
//: {2}(247,319)(295,319){3}
//: {4}(245,317)(245,137)(331,137){5}
//: enddecls

  //: input g8 (Clk) @(120,387) /sn:0 /w:[ 0 ]
  //: supply0 g3 (w11) @(314,184) /sn:0 /w:[ 3 ]
  add g2 (.A(w11), .B(x), .S(PCNext), .CI(!w2), .CO(Cout));   //: @(347,153) /sn:0 /R:1 /w:[ 0 5 1 5 0 ]
  register g1 (.Q(x), .D(PCNew), .EN(w2), .CLR(!Reset), .CK(!Clk));   //: @(184,319) /sn:0 /R:1 /w:[ 0 1 0 1 1 ]
  tran g10(.Z(w2), .I(w11[0]));   //: @(323,167) /sn:0 /R:1 /w:[ 3 2 1 ] /ss:0
  //: input g6 (PCNew) @(122,319) /sn:0 /w:[ 0 ]
  //: input g9 (Reset) @(122,265) /sn:0 /w:[ 0 ]
  //: output g7 (PCNext) @(413,153) /sn:0 /w:[ 0 ]
  //: output g12 (Inst) @(366,317) /sn:0 /w:[ 1 ]
  //: joint g5 (x) @(245, 319) /w:[ 2 4 1 -1 ]
  //: joint g11 (w2) @(214, 153) /w:[ 2 4 1 6 ]
  rom g0 (.A(x), .D(Inst), .OE(w2));   //: @(313,318) /sn:0 /w:[ 3 0 7 ]

endmodule

module ALU(ALUOperation, rt, Zero, ALUResult, rs);
//: interface  /sz:(91, 82) /bd:[ Ti0>ALUOp[3:0](45/91) Ti1>ALUOp[3:0](45/91) Li0>A[31:0](25/82) Li1>B[31:0](51/82) Li2>B[31:0](51/82) Li3>A[31:0](25/82) Bo0<Zero(44/91) Bo1<Zero(44/91) Ro0<ALUResult[31:0](39/82) Ro1<ALUResult[31:0](39/82) ]
output Zero;    //: /sn:0 /dp:1 {0}(295,505)(295,515)(319,515){1}
//: {2}(323,515)(341,515)(341,516)(359,516){3}
//: {4}(321,517)(321,527)(277,527){5}
input [3:0] ALUOperation;    //: /sn:0 /dp:1 {0}(676,331)(676,384)(508,384)(508,479)(65,479){1}
input [31:0] rt;    //: /sn:0 /dp:11 {0}(389,254)(338,254)(338,173){1}
//: {2}(340,171)(399,171){3}
//: {4}(403,171)(418,171){5}
//: {6}(401,173)(401,186)(419,186){7}
//: {8}(336,171)(301,171){9}
//: {10}(297,171)(198,171)(198,170)(100,170){11}
//: {12}(299,173)(299,246){13}
output [31:0] ALUResult;    //: /sn:0 /dp:1 {0}(689,308)(704,308)(704,401){1}
//: {2}(706,403)(768,403){3}
//: {4}(704,405)(704,417)(1084,417)(1084,586)(1064,586){5}
//: {6}(1063,586)(1048,586){7}
//: {8}(1047,586)(1031,586){9}
//: {10}(1030,586)(1015,586){11}
//: {12}(1014,586)(1001,586){13}
//: {14}(1000,586)(986,586){15}
//: {16}(985,586)(970,586){17}
//: {18}(969,586)(954,586){19}
//: {20}(953,586)(937,586){21}
//: {22}(936,586)(920,586){23}
//: {24}(919,586)(908,586){25}
//: {26}(907,586)(890,586){27}
//: {28}(889,586)(874,586){29}
//: {30}(872,586)(857,586){31}
//: {32}(856,586)(838,586){33}
//: {34}(837,586)(823,586){35}
//: {36}(822,586)(806,586){37}
//: {38}(805,586)(791,586){39}
//: {40}(790,586)(776,586){41}
//: {42}(775,586)(760,586){43}
//: {44}(759,586)(743,586){45}
//: {46}(742,586)(730,586){47}
//: {48}(729,586)(714,586){49}
//: {50}(713,586)(707,586)(707,615){51}
//: {52}(707,616)(707,635){53}
//: {54}(707,636)(707,658){55}
//: {56}(707,659)(707,682){57}
//: {58}(707,683)(707,705){59}
//: {60}(707,706)(707,724){61}
//: {62}(707,725)(707,742){63}
//: {64}(707,743)(707,769){65}
//: {66}(707,770)(707,788){67}
//: {68}(707,789)(707,804){69}
supply0 [30:0] w8;    //: /sn:0 {0}(481,371)(502,371)(502,357)(524,357){1}
supply0 [31:0] w49;    //: /sn:0 /dp:1 {0}(660,306)(540,306)(540,308)(530,308){1}
//: {2}(528,306)(528,297){3}
//: {4}(530,295)(660,295){5}
//: {6}(528,293)(528,281){7}
//: {8}(530,279)(538,279)(538,285)(556,285){9}
//: {10}(560,285)(660,285){11}
//: {12}(558,283)(558,281)(660,281){13}
//: {14}(528,277)(528,226){15}
//: {16}(526,295)(516,295)(516,292)(660,292){17}
//: {18}(526,308)(514,308)(514,302)(538,302){19}
//: {20}(542,302)(660,302){21}
//: {22}(540,300)(540,299)(660,299){23}
//: {24}(540,304)(540,314)(555,314)(555,288)(660,288){25}
//: {26}(528,310)(528,342)(533,342){27}
//: {28}(537,342)(552,342){29}
//: {30}(556,342)(562,342)(562,323)(660,323){31}
//: {32}(554,340)(554,320)(660,320){33}
//: {34}(535,340)(535,316)(660,316){35}
supply1 w2;    //: /sn:0 {0}(221,277)(378,277)(378,270)(397,270)(397,280){1}
supply0 w15;    //: /sn:0 {0}(226,201)(403,201)(403,214){1}
input [31:0] rs;    //: /sn:0 /dp:11 {0}(389,222)(326,222){1}
//: {2}(324,220)(324,168){3}
//: {4}(326,166)(391,166){5}
//: {6}(395,166)(418,166){7}
//: {8}(393,168)(393,191)(419,191){9}
//: {10}(322,166)(203,166)(203,155)(83,155){11}
//: {12}(324,224)(324,288)(383,288){13}
wire w16;    //: /sn:0 {0}(484,607)(548,607)(548,770)(702,770){1}
wire w7;    //: /sn:0 {0}(463,575)(390,575)(390,518)(380,518){1}
wire w34;    //: /sn:0 {0}(730,581)(730,562)(484,562){1}
wire w25;    //: /sn:0 {0}(838,581)(838,528)(481,528){1}
wire w4;    //: /sn:0 {0}(1048,581)(1048,463)(481,463){1}
wire w39;    //: /sn:0 /dp:1 {0}(937,581)(937,498)(481,498){1}
wire [31:0] w62;    //: /sn:0 {0}(439,169)(636,169)(636,334)(660,334){1}
wire w36;    //: /sn:0 {0}(702,725)(580,725)(580,597)(484,597){1}
wire w22;    //: /sn:0 {0}(908,581)(908,508)(481,508){1}
wire w3;    //: /sn:0 {0}(1064,581)(1064,458)(481,458){1}
wire w20;    //: /sn:0 {0}(460,496)(390,496)(390,513)(380,513){1}
wire w30;    //: /sn:0 {0}(776,581)(776,547)(484,547){1}
wire w29;    //: /sn:0 {0}(791,581)(791,542)(484,542){1}
wire w42;    //: /sn:0 {0}(397,328)(397,338){1}
wire w37;    //: /sn:0 {0}(702,706)(600,706)(600,592)(484,592){1}
wire [31:0] w18;    //: /sn:0 /dp:1 {0}(418,238)(451,238)(451,232)(612,232)(612,327)(660,327){1}
wire w12;    //: /sn:0 {0}(452,309)(452,367)(524,367){1}
wire [31:0] w10;    //: /sn:0 /dp:1 {0}(412,304)(441,304)(441,305)(451,305){1}
//: {2}(452,305)(578,305)(578,313)(660,313){3}
wire w23;    //: /sn:0 {0}(890,581)(890,513)(481,513){1}
wire [31:0] w63;    //: /sn:0 {0}(440,189)(618,189)(618,330)(660,330){1}
wire w21;    //: /sn:0 {0}(702,743)(566,743)(566,602)(484,602){1}
wire w24;    //: /sn:0 {0}(873,581)(873,518)(481,518){1}
wire w31;    //: /sn:0 {0}(760,581)(760,552)(484,552){1}
wire w32;    //: /sn:0 {0}(743,581)(743,557)(484,557){1}
wire w46;    //: /sn:0 {0}(403,262)(403,272){1}
wire [31:0] w44;    //: /sn:0 {0}(299,262)(299,320)(383,320){1}
wire w27;    //: /sn:0 {0}(823,581)(823,533)(481,533){1}
wire [31:0] w17;    //: /sn:0 /dp:1 {0}(530,362)(607,362)(607,309)(660,309){1}
wire w35;    //: /sn:0 {0}(702,616)(680,616)(680,572)(484,572){1}
wire w33;    //: /sn:0 {0}(714,581)(714,567)(484,567){1}
wire w28;    //: /sn:0 {0}(806,581)(806,537)(484,537){1}
wire w45;    //: /sn:0 /dp:1 {0}(702,659)(641,659)(641,582)(484,582){1}
wire w14;    //: /sn:0 /dp:1 {0}(702,789)(529,789)(529,612)(484,612){1}
wire w11;    //: /sn:0 {0}(1001,581)(1001,478)(481,478){1}
wire w41;    //: /sn:0 /dp:1 {0}(970,581)(970,488)(481,488){1}
wire w47;    //: /sn:0 /dp:1 {0}(702,636)(662,636)(662,577)(484,577){1}
wire w55;    //: /sn:0 {0}(481,483)(986,483)(986,581){1}
wire w5;    //: /sn:0 {0}(1031,581)(1031,468)(481,468){1}
wire w38;    //: /sn:0 /dp:1 {0}(920,581)(920,503)(481,503){1}
wire w43;    //: /sn:0 {0}(702,683)(624,683)(624,587)(484,587){1}
wire w26;    //: /sn:0 {0}(857,581)(857,523)(481,523){1}
wire w9;    //: /sn:0 {0}(1015,581)(1015,473)(481,473){1}
wire w40;    //: /sn:0 /dp:1 {0}(954,581)(954,493)(481,493){1}
//: enddecls

  //: joint g4 (w49) @(535, 342) /w:[ 28 34 27 -1 ]
  tran g44(.Z(w27), .I(ALUResult[16]));   //: @(823,584) /sn:0 /R:1 /w:[ 0 36 35 ] /ss:0
  //: joint g8 (rs) @(393, 166) /w:[ 6 -1 5 8 ]
  //: joint g3 (w49) @(554, 342) /w:[ 30 32 29 -1 ]
  tran g47(.Z(w24), .I(ALUResult[19]));   //: @(873,584) /sn:0 /R:1 /w:[ 0 30 29 ] /ss:0
  //: supply1 g16 (w2) @(221,266) /sn:0 /R:1 /w:[ 0 ]
  concat g17 (.I0(w12), .I1(w8), .Z(w17));   //: @(529,362) /sn:0 /w:[ 1 1 0 ] /dr:0
  //: supply0 g26 (w49) @(528,220) /sn:0 /R:2 /w:[ 15 ]
  //: input g2 (ALUOperation) @(63,479) /sn:0 /w:[ 1 ]
  tran g30(.Z(w21), .I(ALUResult[2]));   //: @(705,743) /sn:0 /R:2 /w:[ 0 64 63 ] /ss:0
  tran g23(.Z(w14), .I(ALUResult[0]));   //: @(705,789) /sn:0 /R:2 /w:[ 0 68 67 ] /ss:0
  nor g24 (.I0(w7), .I1(w20), .Z(Zero));   //: @(369,516) /sn:0 /R:2 /delay:" 2" /w:[ 1 1 3 ]
  tran g39(.Z(w32), .I(ALUResult[11]));   //: @(743,584) /sn:0 /R:1 /w:[ 0 46 45 ] /ss:0
  //: input g1 (rt) @(98,170) /sn:0 /w:[ 11 ]
  tran g29(.Z(w16), .I(ALUResult[1]));   //: @(705,770) /sn:0 /R:2 /w:[ 1 66 65 ] /ss:0
  mux g60 (.I0(w62), .I1(w63), .I2(w18), .I3(w49), .I4(w49), .I5(w49), .I6(w10), .I7(w17), .I8(w49), .I9(w49), .I10(w49), .I11(w49), .I12(w49), .I13(w49), .I14(w49), .I15(w49), .S(ALUOperation), .Z(ALUResult));   //: @(676,308) /sn:0 /R:1 /delay:" 8 8" /w:[ 1 1 1 31 33 35 3 1 0 21 23 5 17 25 11 13 0 0 ] /ss:0 /do:0
  tran g51(.Z(w39), .I(ALUResult[23]));   //: @(937,584) /sn:0 /R:1 /w:[ 0 22 21 ] /ss:0
  tran g18(.Z(w12), .I(w10[31]));   //: @(452,303) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: output g65 (Zero) @(280,527) /sn:0 /R:2 /w:[ 5 ]
  //: joint g25 (rt) @(299, 171) /w:[ 9 -1 10 12 ]
  //: supply0 g10 (w15) @(220,201) /sn:0 /R:3 /w:[ 0 ]
  or g64 (.I0(w14), .I1(w16), .I2(w21), .I3(w36), .I4(w37), .I5(w43), .I6(w45), .I7(w47), .I8(w35), .I9(w33), .I10(w34), .I11(w32), .I12(w31), .I13(w30), .I14(w29), .I15(w28), .Z(w7));   //: @(473,575) /sn:0 /R:2 /delay:" 2" /w:[ 1 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 0 ]
  tran g49(.Z(w22), .I(ALUResult[21]));   //: @(908,584) /sn:0 /R:1 /w:[ 0 26 25 ] /ss:0
  tran g50(.Z(w38), .I(ALUResult[22]));   //: @(920,584) /sn:0 /R:1 /w:[ 0 24 23 ] /ss:0
  or g6 (.I0(rt), .I1(rs), .Z(w63));   //: @(430,189) /sn:0 /w:[ 7 9 0 ]
  //: comment g68 /dolink:0 /link:"" @(147,632) /sn:0
  //: /line:"Set delay to 2x2T and 2T because 32BIT nor gate doesn't work"
  //: /end
  tran g58(.Z(w4), .I(ALUResult[30]));   //: @(1048,584) /sn:0 /R:1 /w:[ 0 8 7 ] /ss:0
  tran g56(.Z(w9), .I(ALUResult[28]));   //: @(1015,584) /sn:0 /R:1 /w:[ 0 12 11 ] /ss:0
  tran g35(.Z(w47), .I(ALUResult[7]));   //: @(705,636) /sn:0 /R:2 /w:[ 0 54 53 ] /ss:0
  //: joint g7 (rt) @(401, 171) /w:[ 4 -1 3 6 ]
  //: joint g22 (w49) @(528, 308) /w:[ 1 2 18 26 ]
  tran g59(.Z(w3), .I(ALUResult[31]));   //: @(1064,584) /sn:0 /R:1 /w:[ 0 6 5 ] /ss:0
  tran g31(.Z(w37), .I(ALUResult[4]));   //: @(705,706) /sn:0 /R:2 /w:[ 0 60 59 ] /ss:0
  led g67 (.I(Zero));   //: @(295,498) /sn:0 /w:[ 0 ] /type:0
  tran g54(.Z(w55), .I(ALUResult[26]));   //: @(986,584) /sn:0 /R:1 /w:[ 1 16 15 ] /ss:0
  tran g45(.Z(w25), .I(ALUResult[17]));   //: @(838,584) /sn:0 /R:1 /w:[ 0 34 33 ] /ss:0
  tran g41(.Z(w30), .I(ALUResult[13]));   //: @(776,584) /sn:0 /R:1 /w:[ 0 42 41 ] /ss:0
  tran g36(.Z(w35), .I(ALUResult[8]));   //: @(705,616) /sn:0 /R:2 /w:[ 0 52 51 ] /ss:0
  tran g33(.Z(w43), .I(ALUResult[5]));   //: @(705,683) /sn:0 /R:2 /w:[ 0 58 57 ] /ss:0
  add g69 (.A(w44), .B(rs), .S(w10), .CI(w2), .CO(w42));   //: @(399,304) /sn:0 /R:1 /w:[ 1 13 0 1 0 ]
  tran g52(.Z(w40), .I(ALUResult[24]));   //: @(954,584) /sn:0 /R:1 /w:[ 0 20 19 ] /ss:0
  tran g42(.Z(w29), .I(ALUResult[14]));   //: @(791,584) /sn:0 /R:1 /w:[ 0 40 39 ] /ss:0
  tran g40(.Z(w31), .I(ALUResult[12]));   //: @(760,584) /sn:0 /R:1 /w:[ 0 44 43 ] /ss:0
  //: joint g66 (Zero) @(321, 515) /w:[ 2 -1 1 4 ]
  //: joint g12 (rs) @(324, 166) /w:[ 4 -1 10 3 ]
  //: joint g28 (w49) @(528, 295) /w:[ 4 6 16 3 ]
  tran g57(.Z(w5), .I(ALUResult[29]));   //: @(1031,584) /sn:0 /R:1 /w:[ 0 10 9 ] /ss:0
  tran g46(.Z(w26), .I(ALUResult[18]));   //: @(857,584) /sn:0 /R:1 /w:[ 0 32 31 ] /ss:0
  tran g34(.Z(w45), .I(ALUResult[6]));   //: @(705,659) /sn:0 /R:2 /w:[ 0 56 55 ] /ss:0
  add g11 (.A(rt), .B(rs), .S(w18), .CI(w15), .CO(w46));   //: @(405,238) /sn:0 /R:1 /w:[ 0 0 0 1 0 ]
  not g14 (.I(rt), .Z(w44));   //: @(299,252) /sn:0 /R:3 /w:[ 13 0 ]
  and g5 (.I0(rs), .I1(rt), .Z(w62));   //: @(429,169) /sn:0 /w:[ 7 5 0 ]
  //: supply0 g19 (w8) @(475,371) /sn:0 /R:3 /w:[ 0 ]
  //: output g21 (ALUResult) @(765,403) /sn:0 /w:[ 3 ]
  //: joint g61 (ALUResult) @(704, 403) /w:[ 2 1 -1 4 ]
  or g20 (.I0(w27), .I1(w25), .I2(w26), .I3(w24), .I4(w23), .I5(w22), .I6(w38), .I7(w39), .I8(w40), .I9(w41), .I10(w55), .I11(w11), .I12(w9), .I13(w5), .I14(w4), .I15(w3), .Z(w20));   //: @(470,496) /sn:0 /R:2 /delay:" 2" /w:[ 1 1 1 1 1 1 1 1 1 1 0 1 1 1 1 1 0 ]
  tran g32(.Z(w36), .I(ALUResult[3]));   //: @(705,725) /sn:0 /R:2 /w:[ 0 62 61 ] /ss:0
  //: joint g63 (w49) @(558, 285) /w:[ 10 12 9 -1 ]
  tran g43(.Z(w28), .I(ALUResult[15]));   //: @(806,584) /sn:0 /R:1 /w:[ 0 38 37 ] /ss:0
  tran g38(.Z(w34), .I(ALUResult[10]));   //: @(730,584) /sn:0 /R:1 /w:[ 0 48 47 ] /ss:0
  //: joint g15 (rs) @(324, 222) /w:[ 1 2 -1 12 ]
  //: input g0 (rs) @(81,155) /sn:0 /w:[ 11 ]
  //: joint g27 (w49) @(540, 302) /w:[ 20 22 19 24 ]
  tran g48(.Z(w23), .I(ALUResult[20]));   //: @(890,584) /sn:0 /R:1 /w:[ 0 28 27 ] /ss:0
  //: joint g62 (w49) @(528, 279) /w:[ 8 14 -1 7 ]
  tran g37(.Z(w33), .I(ALUResult[9]));   //: @(714,584) /sn:0 /R:1 /w:[ 0 50 49 ] /ss:0
  tran g55(.Z(w11), .I(ALUResult[27]));   //: @(1001,584) /sn:0 /R:1 /w:[ 0 14 13 ] /ss:0
  tran g53(.Z(w41), .I(ALUResult[25]));   //: @(970,584) /sn:0 /R:1 /w:[ 0 18 17 ] /ss:0
  //: joint g13 (rt) @(338, 171) /w:[ 2 -1 8 1 ]

endmodule

module EXE(PCNext, ALUResult, Zero, rt, rs, Inm32, BranchTarget, ALUOperation, ALUSrc);
//: interface  /sz:(142, 213) /bd:[ Ti0>ALUOperation[3:0](99/142) Ti1>ALUSrc(36/142) Li0>rt[31:0](114/213) Li1>rs[31:0](81/213) Li2>Inm32[31:0](148/213) Li3>PCNext[31:0](25/213) Ro0<ALUResult[31:0](139/213) Ro1<Zero(57/213) ]
output Zero;    //: /sn:0 {0}(473,294)(333,294){1}
input [31:0] Inm32;    //: /sn:0 {0}(99,165)(119,165){1}
//: {2}(123,165)(283,165){3}
//: {4}(121,167)(121,335)(152,335){5}
input [3:0] ALUOperation;    //: /sn:0 /dp:1 {0}(280,273)(280,230)(96,230){1}
input [31:0] rt;    //: /sn:0 {0}(99,355)(152,355){1}
input ALUSrc;    //: /sn:0 {0}(98,389)(168,389)(168,368){1}
output [31:0] ALUResult;    //: /sn:0 {0}(333,319)(474,319){1}
input [31:0] PCNext;    //: /sn:0 {0}(101,133)(283,133){1}
supply0 CarryIn;    //: /sn:0 /dp:1 {0}(244,85)(297,85)(297,125){1}
output [31:0] BranchTarget;    //: /sn:0 {0}(405,149)(312,149){1}
input [31:0] rs;    //: /sn:0 {0}(98,302)(235,302){1}
wire [31:0] w4;    //: /sn:0 /dp:1 {0}(181,345)(235,345){1}
wire Overflow;    //: /sn:0 /dp:1 {0}(297,173)(297,199)(351,199){1}
//: enddecls

  //: input g8 (PCNext) @(99,133) /sn:0 /w:[ 0 ]
  //: output g4 (ALUResult) @(471,319) /sn:0 /w:[ 1 ]
  //: output g3 (Zero) @(470,294) /sn:0 /w:[ 0 ]
  //: input g2 (rt) @(97,355) /sn:0 /w:[ 0 ]
  //: input g1 (rs) @(96,302) /sn:0 /w:[ 0 ]
  //: supply0 g10 (CarryIn) @(238,85) /sn:0 /R:3 /w:[ 0 ]
  add g6 (.A(Inm32), .B(PCNext), .S(BranchTarget), .CI(CarryIn), .CO(Overflow));   //: @(299,149) /sn:0 /R:1 /w:[ 3 1 1 1 0 ]
  //: input g7 (Inm32) @(97,165) /sn:0 /w:[ 0 ]
  //: output g9 (BranchTarget) @(402,149) /sn:0 /w:[ 0 ]
  //: joint g12 (Inm32) @(121, 165) /w:[ 2 -1 1 4 ]
  mux g11 (.I0(rt), .I1(Inm32), .S(ALUSrc), .Z(w4));   //: @(168,345) /sn:0 /R:1 /w:[ 1 5 1 0 ] /ss:0 /do:0
  //: input g5 (ALUOperation) @(94,230) /sn:0 /w:[ 1 ]
  ALU g0 (.ALUOperation(ALUOperation), .rt(w4), .rs(rs), .Zero(Zero), .ALUResult(ALUResult));   //: @(236, 274) /sz:(96, 97) /sn:0 /p:[ Ti0>0 Li0>1 Li1>1 Ro0<1 Ro1<0 ]
  //: input g13 (ALUSrc) @(96,389) /sn:0 /w:[ 0 ]

endmodule

module BRegs32x32(Read2, Write, Read1, Data2, Data1, clr, clk, RegWrite, WriteData);
//: interface  /sz:(147, 182) /bd:[ Ti0>clr(66/147) Ti1>clr(66/147) Ti2>clr(66/147) Ti3>clr(66/147) Ti4>clr(66/147) Ti5>clr(66/147) Ti6>clr(66/147) Ti7>clr(66/147) Ti8>clr(66/147) Li0>WriteData[31:0](148/182) Li1>Write[4:0](108/182) Li2>Read2[4:0](72/182) Li3>Read1[4:0](32/182) Li4>Read1[4:0](32/182) Li5>Read2[4:0](72/182) Li6>Write[4:0](108/182) Li7>WriteData[31:0](148/182) Li8>WriteData[31:0](148/182) Li9>Write[4:0](108/182) Li10>Read2[4:0](72/182) Li11>Read1[4:0](32/182) Li12>WriteData[31:0](148/182) Li13>Write[4:0](108/182) Li14>Read2[4:0](72/182) Li15>Read1[4:0](32/182) Li16>Read1[4:0](32/182) Li17>Read2[4:0](72/182) Li18>Write[4:0](108/182) Li19>WriteData[31:0](148/182) Li20>WriteData[31:0](148/182) Li21>Write[4:0](108/182) Li22>Read2[4:0](72/182) Li23>Read1[4:0](32/182) Li24>WriteData[31:0](148/182) Li25>Write[4:0](108/182) Li26>Read2[4:0](72/182) Li27>Read1[4:0](32/182) Li28>Read1[4:0](32/182) Li29>Read2[4:0](72/182) Li30>Write[4:0](108/182) Li31>WriteData[31:0](148/182) Li32>WriteData[31:0](148/182) Li33>Write[4:0](108/182) Li34>Read2[4:0](72/182) Li35>Read1[4:0](32/182) Bi0>RegWrite(40/147) Bi1>clk(108/147) Bi2>clk(108/147) Bi3>RegWrite(40/147) Bi4>RegWrite(40/147) Bi5>clk(108/147) Bi6>RegWrite(40/147) Bi7>clk(108/147) Bi8>clk(108/147) Bi9>RegWrite(40/147) Bi10>RegWrite(40/147) Bi11>clk(108/147) Bi12>RegWrite(40/147) Bi13>clk(108/147) Bi14>clk(108/147) Bi15>RegWrite(40/147) Bi16>RegWrite(40/147) Bi17>clk(108/147) Ro0<Data2[31:0](139/182) Ro1<Data1[31:0](47/182) Ro2<Data1[31:0](47/182) Ro3<Data2[31:0](139/182) Ro4<Data2[31:0](139/182) Ro5<Data1[31:0](47/182) Ro6<Data2[31:0](139/182) Ro7<Data1[31:0](47/182) Ro8<Data1[31:0](47/182) Ro9<Data2[31:0](139/182) Ro10<Data2[31:0](139/182) Ro11<Data1[31:0](47/182) Ro12<Data2[31:0](139/182) Ro13<Data1[31:0](47/182) Ro14<Data1[31:0](47/182) Ro15<Data2[31:0](139/182) Ro16<Data2[31:0](139/182) Ro17<Data1[31:0](47/182) ]
output [31:0] Data2;    //: /sn:0 {0}(668,485)(668,472)(669,472)(669,445){1}
input [4:0] Write;    //: /sn:0 {0}(-238,-38)(-138,-38)(-138,-37)(-66,-37){1}
//: {2}(-65,-37)(-28,-37){3}
//: {4}(-27,-37)(-16,-37){5}
input [31:0] WriteData;    //: /sn:0 {0}(669,157)(669,75)(481,75){1}
//: {2}(477,75)(292,75){3}
//: {4}(288,75)(89,75){5}
//: {6}(85,75)(-104,75)(-104,73)(-237,73){7}
//: {8}(87,77)(87,157){9}
//: {10}(290,77)(290,107)(291,107)(291,152){11}
//: {12}(479,77)(479,157){13}
supply1 w21;    //: /sn:0 {0}(82,3)(57,3)(57,-11){1}
output [31:0] Data1;    //: /sn:0 {0}(59,382)(59,465){1}
input RegWrite;    //: /sn:0 {0}(-237,263)(-71,263){1}
//: {2}(-67,263)(171,263){3}
//: {4}(175,263)(370,263){5}
//: {6}(374,263)(552,263)(552,219)(556,219){7}
//: {8}(372,261)(372,219)(383,219){9}
//: {10}(173,261)(173,214)(183,214){11}
//: {12}(-69,261)(-69,219)(-38,219){13}
input clr;    //: /sn:0 {0}(721,193)(731,193)(731,-83)(543,-83){1}
//: {2}(539,-83)(355,-83){3}
//: {4}(351,-83)(150,-83){5}
//: {6}(146,-83)(-44,-83)(-44,-92)(-235,-92){7}
//: {8}(148,-81)(148,193)(139,193){9}
//: {10}(353,-81)(353,188)(343,188){11}
//: {12}(541,-81)(541,193)(531,193){13}
input clk;    //: /sn:0 {0}(556,214)(542,214)(542,285)(364,285){1}
//: {2}(362,283)(362,214)(383,214){3}
//: {4}(360,285)(167,285){5}
//: {6}(165,283)(165,209)(183,209){7}
//: {8}(163,285)(-56,285){9}
//: {10}(-58,283)(-58,214)(-38,214){11}
//: {12}(-60,285)(-237,285){13}
input [4:0] Read1;    //: {0}(-237,96)(-208,96)(-208,95)(-124,95){1}
//: {2}(-123,95)(-96,95){3}
//: {4}(-95,95)(-78,95){5}
input [4:0] Read2;    //: {0}(-237,145)(-141,145){1}
//: {2}(-140,145)(-123,145)(-123,144)(-94,144){3}
//: {4}(-93,144)(-79,144){5}
wire w16;    //: /sn:0 {0}(39,205)(-50,205)(-50,39)(88,39)(88,19){1}
wire [1:0] w6;    //: /sn:0 {0}(36,369)(-123,369)(-123,99){1}
wire w4;    //: /sn:0 {0}(112,19)(112,46)(370,46)(370,205)(431,205){1}
wire w22;    //: /sn:0 {0}(404,217)(431,217){1}
wire [31:0] w0;    //: /sn:0 {0}(651,416)(651,398)(105,398)(105,228){1}
wire [31:0] R2;    //: {0}(65,353)(65,319)(469,319)(469,228){1}
wire [31:0] w3;    //: /sn:0 {0}(77,353)(77,334)(659,334)(659,228){1}
wire w20;    //: /sn:0 {0}(124,19)(124,29)(556,29)(556,205)(621,205){1}
wire [2:0] w18;    //: /sn:0 {0}(431,180)(402,180)(402,125){1}
//: {2}(404,123)(589,123)(589,180)(621,180){3}
//: {4}(400,123)(279,123)(279,122)(212,122){5}
//: {6}(208,122)(8,122){7}
//: {8}(4,122)(-93,122)(-93,139){9}
//: {10}(6,124)(6,180)(39,180){11}
//: {12}(210,124)(210,175)(243,175){13}
wire [2:0] w19;    //: /sn:0 {0}(431,169)(419,169)(419,109){1}
//: {2}(421,107)(606,107)(606,169)(621,169){3}
//: {4}(417,107)(297,107)(297,106)(231,106){5}
//: {6}(227,106)(25,106){7}
//: {8}(21,106)(-95,106)(-95,99){9}
//: {10}(23,108)(23,169)(39,169){11}
//: {12}(229,108)(229,164)(243,164){13}
wire [1:0] w10;    //: /sn:0 {0}(-140,149)(-140,432)(646,432){1}
wire w23;    //: /sn:0 {0}(577,217)(621,217){1}
wire [2:0] w24;    //: /sn:0 {0}(431,193)(381,193)(381,141){1}
//: {2}(383,139)(568,139)(568,193)(621,193){3}
//: {4}(379,139)(260,139)(260,138)(195,138){5}
//: {6}(191,138)(-13,138){7}
//: {8}(-17,138)(-65,138)(-65,-33){9}
//: {10}(-15,140)(-15,193)(39,193){11}
//: {12}(193,140)(193,188)(243,188){13}
wire w1;    //: /sn:0 {0}(-17,217)(39,217){1}
wire w31;    //: /sn:0 {0}(243,200)(178,200)(178,60)(100,60)(100,19){1}
wire [31:0] R3;    //: {0}(687,228)(687,416){1}
wire [31:0] R1;    //: {0}(281,223)(281,308)(53,308)(53,353){1}
wire w2;    //: /sn:0 {0}(243,212)(204,212){1}
wire [1:0] w11;    //: /sn:0 {0}(-27,-33)(-27,-23)(106,-23)(106,-10){1}
wire [31:0] R0;    //: {0}(77,228)(77,299)(41,299)(41,353){1}
wire [31:0] w5;    //: /sn:0 {0}(675,416)(675,372)(497,372)(497,228){1}
wire [31:0] w9;    //: /sn:0 {0}(663,416)(663,387)(309,387)(309,223){1}
//: enddecls

  //: joint g44 (clr) @(353, -83) /w:[ 3 -1 4 10 ]
  //: input g4 (Read2) @(-239,145) /sn:0 /w:[ 0 ]
  //: joint g8 (w18) @(6, 122) /w:[ 7 -1 8 10 ]
  //: joint g47 (clr) @(541, -83) /w:[ 1 -1 2 12 ]
  //: joint g16 (clk) @(165, 285) /w:[ 5 6 8 -1 ]
  //: input g3 (Write) @(-240,-38) /sn:0 /w:[ 0 ]
  //: joint g26 (w19) @(229, 106) /w:[ 5 -1 6 12 ]
  //: input g17 (Read1) @(-239,96) /sn:0 /w:[ 0 ]
  //: output g2 (Data2) @(668,482) /sn:0 /R:3 /w:[ 0 ]
  tran g30(.Z(w10), .I(Read2[4:3]));   //: @(-140,143) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  tran g23(.Z(w24), .I(Write[2:0]));   //: @(-65,-39) /sn:0 /R:1 /w:[ 9 1 2 ] /ss:1
  Regs8x32 g24 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w31), .clk(w2), .clr(clr), .AOUT(R1), .BOUT(w9));   //: @(244, 153) /sz:(98, 69) /sn:0 /p:[ Ti0>11 Li0>13 Li1>13 Li2>13 Li3>0 Li4>0 Ri0>11 Bo0<0 Bo1<1 ]
  //: joint g39 (RegWrite) @(372, 263) /w:[ 6 8 5 -1 ]
  //: output g1 (Data1) @(59,462) /sn:0 /R:3 /w:[ 1 ]
  Regs8x32 g29 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w4), .clk(w22), .clr(clr), .AOUT(R2), .BOUT(w5));   //: @(432, 158) /sz:(98, 69) /sn:0 /p:[ Ti0>13 Li0>0 Li1>0 Li2>0 Li3>1 Li4>1 Ri0>13 Bo0<1 Bo1<1 ]
  //: comment g51 /dolink:0 /link:"" @(395,229) /sn:0
  //: /line:"Regs 16-23"
  //: /end
  tran g18(.Z(w19), .I(Read1[2:0]));   //: @(-95,93) /sn:0 /R:1 /w:[ 9 3 4 ] /ss:1
  //: joint g25 (w18) @(210, 122) /w:[ 5 -1 6 12 ]
  //: supply1 g10 (w21) @(68,-11) /sn:0 /w:[ 1 ]
  //: comment g49 /dolink:0 /link:"" @(210,225) /sn:0
  //: /line:"Regs 8-15"
  //: /end
  Regs8x32 g6 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w16), .clk(w1), .clr(clr), .AOUT(R0), .BOUT(w0));   //: @(40, 158) /sz:(98, 69) /sn:0 /p:[ Ti0>9 Li0>11 Li1>11 Li2>11 Li3>0 Li4>1 Ri0>9 Bo0<0 Bo1<1 ]
  //: comment g50 /dolink:0 /link:"" @(585,229) /sn:0
  //: /line:"Regs 24-31"
  //: /end
  and g35 (.I0(clk), .I1(RegWrite), .Z(w22));   //: @(394,217) /sn:0 /delay:" 1" /w:[ 3 9 0 ]
  demux g9 (.I(w11), .E(w21), .Z0(w16), .Z1(w31), .Z2(w4), .Z3(w20));   //: @(106,3) /sn:0 /w:[ 1 0 1 1 0 0 ]
  //: joint g7 (w19) @(23, 106) /w:[ 7 -1 8 10 ]
  tran g22(.Z(w18), .I(Read2[2:0]));   //: @(-93,142) /sn:0 /R:1 /w:[ 9 3 4 ] /ss:0
  tran g31(.Z(w6), .I(Read1[4:3]));   //: @(-123,93) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  and g33 (.I0(clk), .I1(RegWrite), .Z(w1));   //: @(-27,217) /sn:0 /delay:" 1" /w:[ 11 13 0 ]
  //: joint g45 (WriteData) @(479, 75) /w:[ 1 -1 2 12 ]
  //: joint g41 (w19) @(419, 107) /w:[ 2 -1 4 1 ]
  and g36 (.I0(clk), .I1(RegWrite), .Z(w23));   //: @(567,217) /sn:0 /delay:" 1" /w:[ 0 7 0 ]
  //: joint g40 (w18) @(402, 123) /w:[ 2 -1 4 1 ]
  //: input g42 (clr) @(-237,-92) /sn:0 /w:[ 7 ]
  //: input g12 (clk) @(-239,285) /sn:0 /w:[ 13 ]
  Regs8x32 g46 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w20), .clk(w23), .clr(clr), .AOUT(w3), .BOUT(R3));   //: @(622, 158) /sz:(98, 69) /sn:0 /p:[ Ti0>0 Li0>3 Li1>3 Li2>3 Li3>1 Li4>1 Ri0>0 Bo0<1 Bo1<0 ]
  //: joint g28 (w24) @(381, 139) /w:[ 2 -1 4 1 ]
  and g34 (.I0(clk), .I1(RegWrite), .Z(w2));   //: @(194,212) /sn:0 /delay:" 1" /w:[ 7 11 1 ]
  tran g5(.Z(w11), .I(Write[4:3]));   //: @(-27,-39) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  mux g14 (.I0(R0), .I1(R1), .I2(R2), .I3(w3), .S(w6), .Z(Data1));   //: @(59,369) /sn:0 /w:[ 1 1 0 0 0 0 ] /ss:0 /do:0
  //: joint g11 (w24) @(-15, 138) /w:[ 7 -1 8 10 ]
  //: joint g21 (w24) @(193, 138) /w:[ 5 -1 6 12 ]
  //: joint g19 (clk) @(-58, 285) /w:[ 9 10 12 -1 ]
  //: joint g20 (WriteData) @(87, 75) /w:[ 5 -1 6 8 ]
  //: input g32 (RegWrite) @(-239,263) /sn:0 /w:[ 0 ]
  //: input g0 (WriteData) @(-239,73) /sn:0 /w:[ 7 ]
  //: joint g43 (clr) @(148, -83) /w:[ 5 -1 6 8 ]
  //: joint g15 (clk) @(362, 285) /w:[ 1 2 4 -1 ]
  //: joint g38 (RegWrite) @(173, 263) /w:[ 4 10 3 -1 ]
  //: comment g48 /dolink:0 /link:"" @(11,228) /sn:0
  //: /line:"Regs 0-7"
  //: /end
  //: joint g27 (WriteData) @(290, 75) /w:[ 3 -1 4 10 ]
  //: joint g37 (RegWrite) @(-69, 263) /w:[ 2 12 1 -1 ]
  mux g13 (.I0(w0), .I1(w9), .I2(w5), .I3(R3), .S(w10), .Z(Data2));   //: @(669,432) /sn:0 /w:[ 0 0 0 1 1 1 ] /ss:0 /do:0

endmodule

module Regs8x32(SB, SA, BOUT, AOUT, clr, clk, RegWr, SD, DIN);
//: interface  /sz:(98, 69) /bd:[ Ti0>DIN[31:0](47/98) Ti1>DIN[31:0](47/98) Ti2>DIN[31:0](47/98) Ti3>DIN[31:0](47/98) Ti4>DIN[31:0](47/98) Ti5>DIN[31:0](47/98) Ti6>DIN[31:0](47/98) Ti7>DIN[31:0](47/98) Ti8>DIN[31:0](47/98) Li0>SD[2:0](35/69) Li1>SA[2:0](11/69) Li2>SB[2:0](22/69) Li3>RegWr(47/69) Li4>clk(59/69) Li5>clk(59/69) Li6>RegWr(47/69) Li7>SB[2:0](22/69) Li8>SA[2:0](11/69) Li9>SD[2:0](35/69) Li10>SD[2:0](35/69) Li11>SA[2:0](11/69) Li12>SB[2:0](22/69) Li13>RegWr(47/69) Li14>clk(59/69) Li15>SD[2:0](35/69) Li16>SA[2:0](11/69) Li17>SB[2:0](22/69) Li18>RegWr(47/69) Li19>clk(59/69) Li20>clk(59/69) Li21>RegWr(47/69) Li22>SB[2:0](22/69) Li23>SA[2:0](11/69) Li24>SD[2:0](35/69) Li25>SD[2:0](35/69) Li26>SA[2:0](11/69) Li27>SB[2:0](22/69) Li28>RegWr(47/69) Li29>clk(59/69) Li30>SD[2:0](35/69) Li31>SA[2:0](11/69) Li32>SB[2:0](22/69) Li33>RegWr(47/69) Li34>clk(59/69) Li35>clk(59/69) Li36>RegWr(47/69) Li37>SB[2:0](22/69) Li38>SA[2:0](11/69) Li39>SD[2:0](35/69) Li40>SD[2:0](35/69) Li41>SA[2:0](11/69) Li42>SB[2:0](22/69) Li43>RegWr(47/69) Li44>clk(59/69) Ri0>clr(35/69) Ri1>clr(35/69) Ri2>clr(35/69) Ri3>clr(35/69) Ri4>clr(35/69) Ri5>clr(35/69) Ri6>clr(35/69) Ri7>clr(35/69) Ri8>clr(35/69) Bo0<AOUT[31:0](37/98) Bo1<BOUT[31:0](65/98) Bo2<BOUT[31:0](65/98) Bo3<AOUT[31:0](37/98) Bo4<AOUT[31:0](37/98) Bo5<BOUT[31:0](65/98) Bo6<AOUT[31:0](37/98) Bo7<BOUT[31:0](65/98) Bo8<BOUT[31:0](65/98) Bo9<AOUT[31:0](37/98) Bo10<AOUT[31:0](37/98) Bo11<BOUT[31:0](65/98) Bo12<AOUT[31:0](37/98) Bo13<BOUT[31:0](65/98) Bo14<BOUT[31:0](65/98) Bo15<AOUT[31:0](37/98) Bo16<AOUT[31:0](37/98) Bo17<BOUT[31:0](65/98) ]
input [31:0] DIN;    //: /sn:0 {0}(531,269)(531,318){1}
//: {2}(533,320)(627,320){3}
//: {4}(631,320)(715,320){5}
//: {6}(719,320)(807,320)(807,429){7}
//: {8}(717,322)(717,352){9}
//: {10}(629,322)(629,433){11}
//: {12}(529,320)(435,320){13}
//: {14}(431,320)(342,320){15}
//: {16}(338,320)(264,320){17}
//: {18}(260,320)(181,320)(181,352){19}
//: {20}(262,322)(262,439){21}
//: {22}(340,322)(340,351){23}
//: {24}(433,322)(433,436){25}
//: {26}(531,322)(531,348){27}
output [31:0] BOUT;    //: /sn:0 {0}(516,697)(516,672){1}
input [2:0] SD;    //: /sn:0 {0}(782,138)(852,138)(852,156){1}
input [2:0] SB;    //: /sn:0 {0}(466,659)(493,659){1}
supply1 w21;    //: /sn:0 {0}(828,169)(801,169)(801,153){1}
input RegWr;    //: /sn:0 {0}(48,363)(68,363)(68,378)(82,378){1}
input clr;    //: /sn:0 /dp:1 {0}(959,337)(1032,337){1}
input [2:0] SA;    //: /sn:0 {0}(256,657)(231,657){1}
input clk;    //: /sn:0 {0}(82,383)(68,383)(68,398)(55,398){1}
output [31:0] AOUT;    //: /sn:0 {0}(279,670)(279,702){1}
wire [31:0] w16;    //: /sn:0 {0}(531,369)(531,574)(520,574){1}
//: {2}(516,574)(282,574)(282,641){3}
//: {4}(518,576)(518,587)(519,587)(519,643){5}
wire w7;    //: /sn:0 {0}(472,451)(513,451)(513,405)(848,405)(848,185){1}
wire [31:0] R5;    //: {0}(288,641)(288,586)(525,586){1}
//: {2}(529,586)(629,586)(629,454){3}
//: {4}(527,588)(527,617)(525,617)(525,643){5}
wire w4;    //: /sn:0 {0}(943,337)(906,337){1}
//: {2}(902,337)(767,337){3}
//: {4}(763,337)(588,337){5}
//: {6}(584,337)(390,337){7}
//: {8}(386,337)(231,337)(231,357)(220,357){9}
//: {10}(388,339)(388,356)(379,356){11}
//: {12}(586,339)(586,353)(570,353){13}
//: {14}(765,339)(765,357)(756,357){15}
//: {16}(904,339)(904,417)(865,417){17}
//: {18}(861,417)(675,417){19}
//: {20}(671,417)(489,417){21}
//: {22}(485,417)(302,417)(302,444)(301,444){23}
//: {24}(487,419)(487,441)(472,441){25}
//: {26}(673,419)(673,438)(668,438){27}
//: {28}(863,419)(863,434)(846,434){29}
wire w3;    //: /sn:0 {0}(835,185)(835,397)(330,397)(330,454)(301,454){1}
wire w0;    //: /sn:0 {0}(770,439)(764,439)(764,481)(579,481){1}
//: {2}(577,479)(577,443)(592,443){3}
//: {4}(575,481)(390,481){5}
//: {6}(388,479)(388,446)(396,446){7}
//: {8}(386,481)(214,481){9}
//: {10}(212,479)(212,449)(225,449){11}
//: {12}(210,481)(125,481)(125,383){13}
//: {14}(127,381)(291,381){15}
//: {16}(295,381)(477,381){17}
//: {18}(481,381)(660,381)(660,362)(680,362){19}
//: {20}(479,379)(479,358)(494,358){21}
//: {22}(293,379)(293,361)(303,361){23}
//: {24}(125,379)(125,362)(144,362){25}
//: {26}(123,381)(103,381){27}
wire [31:0] R2;    //: {0}(262,641)(262,537){1}
//: {2}(264,535)(499,535)(499,643){3}
//: {4}(262,533)(262,460){5}
wire [31:0] R7;    //: {0}(807,450)(807,609)(541,609){1}
//: {2}(537,609)(302,609)(302,641){3}
//: {4}(539,611)(539,643){5}
wire w12;    //: /sn:0 {0}(756,367)(787,367)(787,258)(868,258)(868,185){1}
wire w10;    //: /sn:0 {0}(846,444)(875,444)(875,185){1}
wire [31:0] R4;    //: {0}(340,372)(340,545){1}
//: {2}(342,547)(505,547)(505,643){3}
//: {4}(338,547)(268,547)(268,641){5}
wire [31:0] R3;    //: {0}(512,643)(512,559)(435,559){1}
//: {2}(433,557)(433,457){3}
//: {4}(431,559)(275,559)(275,641){5}
wire w8;    //: /sn:0 {0}(220,367)(249,367)(249,213)(828,213)(828,185){1}
wire Z5;    //: /sn:0 {0}(861,185)(861,413)(700,413)(700,448)(668,448){1}
wire w14;    //: /sn:0 {0}(379,366)(414,366)(414,229)(841,229)(841,185){1}
wire [31:0] R0;    //: {0}(492,643)(492,523)(257,523){1}
//: {2}(253,523)(181,523)(181,373){3}
//: {4}(255,525)(255,641){5}
wire w15;    //: /sn:0 {0}(570,363)(608,363)(608,244)(855,244)(855,185){1}
wire [31:0] R10;    //: /sn:0 {0}(295,641)(295,600)(530,600){1}
//: {2}(534,600)(717,600)(717,373){3}
//: {4}(532,602)(532,643){5}
//: enddecls

  //: input g4 (SB) @(464,659) /sn:0 /w:[ 0 ]
  //: joint g8 (w16) @(518, 574) /w:[ 1 -1 2 4 ]
  //: joint g16 (R3) @(433, 559) /w:[ 1 2 4 -1 ]
  //: input g3 (SA) @(229,657) /sn:0 /w:[ 1 ]
  //: joint g26 (DIN) @(340, 320) /w:[ 15 -1 16 22 ]
  //: joint g17 (R4) @(340, 547) /w:[ 2 1 4 -1 ]
  //: output g2 (BOUT) @(516,694) /sn:0 /R:3 /w:[ 0 ]
  register R5 (.Q(R5), .D(DIN), .EN(Z5), .CLR(w4), .CK(!w0));   //: @(629,443) /w:[ 3 11 1 27 3 ]
  //: joint g30 (w0) @(212, 481) /w:[ 9 10 12 -1 ]
  //: joint g23 (w4) @(765, 337) /w:[ 3 -1 4 14 ]
  //: joint g24 (DIN) @(531, 320) /w:[ 2 1 12 26 ]
  //: joint g39 (DIN) @(262, 320) /w:[ 17 -1 18 20 ]
  //: output g1 (AOUT) @(279,699) /sn:0 /R:3 /w:[ 1 ]
  //: joint g29 (w0) @(388, 481) /w:[ 5 6 8 -1 ]
  register R2 (.Q(R4), .D(DIN), .EN(w14), .CLR(w4), .CK(!w0));   //: @(340,361) /w:[ 0 23 0 11 23 ]
  //: joint g18 (R2) @(262, 535) /w:[ 2 4 -1 1 ]
  register R7 (.Q(R7), .D(DIN), .EN(w10), .CLR(w4), .CK(!w0));   //: @(807,439) /w:[ 0 7 0 29 0 ]
  not g25 (.I(clr), .Z(w4));   //: @(953,337) /sn:0 /R:2 /w:[ 0 0 ]
  //: supply1 g10 (w21) @(812,153) /sn:0 /w:[ 1 ]
  register R6 (.Q(R10), .D(DIN), .EN(w12), .CLR(w4), .CK(!w0));   //: @(717,362) /w:[ 3 9 0 15 19 ]
  //: joint g6 (R7) @(539, 609) /w:[ 1 -1 2 4 ]
  and g35 (.I0(RegWr), .I1(clk), .Z(w0));   //: @(93,381) /sn:0 /delay:" 1" /w:[ 1 0 27 ]
  demux g9 (.I(SD), .E(w21), .Z0(!w8), .Z1(!w3), .Z2(!w14), .Z3(!w7), .Z4(!w15), .Z5(!Z5), .Z6(!w12), .Z7(!w10));   //: @(852,169) /sn:0 /w:[ 1 0 1 0 1 1 1 0 1 1 ]
  register R4 (.Q(w16), .D(DIN), .EN(w15), .CLR(w4), .CK(!w0));   //: @(531,358) /w:[ 0 27 0 13 21 ]
  //: joint g7 (R10) @(532, 600) /w:[ 2 -1 1 4 ]
  //: joint g22 (w4) @(586, 337) /w:[ 5 -1 6 12 ]
  //: joint g31 (w4) @(863, 417) /w:[ 17 -1 18 28 ]
  register R1 (.Q(R2), .D(DIN), .EN(w3), .CLR(w4), .CK(!w0));   //: @(262,449) /w:[ 5 21 1 23 11 ]
  register R3 (.Q(R3), .D(DIN), .EN(w7), .CLR(w4), .CK(!w0));   //: @(433,446) /w:[ 3 25 0 25 7 ]
  //: joint g33 (w4) @(673, 417) /w:[ 19 -1 20 26 ]
  //: joint g41 (DIN) @(717, 320) /w:[ 6 -1 5 8 ]
  //: joint g36 (w4) @(904, 337) /w:[ 1 -1 2 16 ]
  //: joint g40 (DIN) @(433, 320) /w:[ 13 -1 14 24 ]
  //: joint g42 (DIN) @(629, 320) /w:[ 4 -1 3 10 ]
  //: joint g12 (w0) @(479, 381) /w:[ 18 20 17 -1 ]
  //: input g28 (clr) @(1034,337) /sn:0 /R:2 /w:[ 1 ]
  //: input g34 (clk) @(53,398) /sn:0 /w:[ 1 ]
  mux g14 (.I0(R0), .I1(R2), .I2(R4), .I3(R3), .I4(w16), .I5(R5), .I6(R10), .I7(R7), .S(SA), .Z(AOUT));   //: @(279,657) /sn:0 /w:[ 5 0 5 5 3 0 0 3 0 0 ] /ss:0 /do:0
  //: input g5 (RegWr) @(46,363) /sn:0 /w:[ 0 ]
  //: joint g11 (w0) @(293, 381) /w:[ 16 22 15 -1 ]
  //: joint g21 (w4) @(388, 337) /w:[ 7 -1 8 10 ]
  //: joint g19 (R0) @(255, 523) /w:[ 1 -1 2 4 ]
  //: input g20 (SD) @(780,138) /sn:0 /w:[ 0 ]
  //: joint g32 (w4) @(487, 417) /w:[ 21 -1 22 24 ]
  register R0 (.Q(R0), .D(DIN), .EN(w8), .CLR(w4), .CK(!w0));   //: @(181,362) /w:[ 3 19 0 9 25 ]
  //: input g0 (DIN) @(531,267) /sn:0 /R:3 /w:[ 0 ]
  //: joint g15 (R5) @(527, 586) /w:[ 2 -1 1 4 ]
  //: joint g38 (w0) @(577, 481) /w:[ 1 2 4 -1 ]
  //: joint g27 (w0) @(125, 381) /w:[ 14 24 26 13 ]
  mux g13 (.I0(R0), .I1(R2), .I2(R4), .I3(R3), .I4(w16), .I5(R5), .I6(R10), .I7(R7), .S(SB), .Z(BOUT));   //: @(516,659) /sn:0 /w:[ 0 3 3 0 5 5 5 5 1 1 ] /ss:0 /do:0

endmodule

module Read(clk, Inm32, Inst, rs, RegDst, WriteData, clr, rt, RegWrite);
//: interface  /sz:(166, 219) /bd:[ Ti0>RegWrite(84/166) Li0>Inst[31:0](30/219) Li1>RegDst(121/219) Bi0>WriteData[31:0](40/166) Bi1>clr(123/166) Bi2>clk(93/166) Ro0<rs[31:0](51/219) Ro1<rt[31:0](92/219) Ro2<Inm32[31:0](141/219) ]
output [31:0] Inm32;    //: /sn:0 /dp:1 {0}(484,464)(614,464){1}
input [31:0] WriteData;    //: /sn:0 /dp:1 {0}(389,297)(365,297)(365,319)(145,319){1}
output [31:0] rt;    //: /sn:0 /dp:1 {0}(538,288)(627,288){1}
input [31:0] Inst;    //: /sn:0 {0}(212,308)(212,298){1}
//: {2}(212,297)(212,268){3}
//: {4}(212,267)(212,221){5}
//: {6}(212,220)(212,181){7}
//: {8}(212,180)(212,138){9}
input RegDst;    //: /sn:0 {0}(146,348)(318,348)(318,281){1}
input clr;    //: /sn:0 {0}(406,77)(462,77)(462,148){1}
input RegWrite;    //: /sn:0 {0}(145,375)(430,375)(430,332){1}
input clk;    //: /sn:0 {0}(144,397)(498,397)(498,332){1}
output [31:0] rs;    //: /sn:0 {0}(622,196)(538,196){1}
wire [4:0] w6;    //: /sn:0 {0}(216,268)(302,268){1}
wire [4:0] w3;    //: /sn:0 {0}(216,181)(389,181){1}
wire [4:0] w0;    //: /sn:0 {0}(302,248)(262,248)(262,223){1}
//: {2}(264,221)(389,221){3}
//: {4}(260,221)(216,221){5}
wire [4:0] w10;    //: /sn:0 {0}(331,258)(389,258){1}
wire [15:0] w8;    //: /sn:0 /dp:1 {0}(442,462)(224,462)(224,298)(216,298){1}
//: enddecls

  //: joint g4 (w0) @(262, 221) /w:[ 2 -1 4 1 ]
  //: input g8 (clk) @(142,397) /sn:0 /w:[ 0 ]
  mux g3 (.I0(w0), .I1(w6), .S(RegDst), .Z(w10));   //: @(318,258) /sn:0 /R:1 /w:[ 0 1 1 0 ] /ss:0 /do:1
  //: output g16 (Inm32) @(611,464) /sn:0 /w:[ 1 ]
  //: input g17 (Inst) @(212,136) /sn:0 /R:3 /w:[ 9 ]
  tran g2(.Z(w0), .I(Inst[20:16]));   //: @(210,221) /sn:0 /R:2 /w:[ 5 5 6 ] /ss:1
  tran g1(.Z(w3), .I(Inst[25:21]));   //: @(210,181) /sn:0 /R:2 /w:[ 0 7 8 ] /ss:1
  //: output g10 (rs) @(619,196) /sn:0 /w:[ 0 ]
  //: input g6 (RegDst) @(144,348) /sn:0 /w:[ 0 ]
  //: input g7 (WriteData) @(143,319) /sn:0 /w:[ 1 ]
  //: input g9 (clr) @(404,77) /sn:0 /w:[ 0 ]
  tran g14(.Z(w8), .I(Inst[15:0]));   //: @(210,298) /sn:0 /R:2 /w:[ 1 1 2 ] /ss:1
  tran g5(.Z(w6), .I(Inst[15:11]));   //: @(210,268) /sn:0 /R:2 /w:[ 0 3 4 ] /ss:1
  //: output g11 (rt) @(624,288) /sn:0 /w:[ 1 ]
  BRegs32x32 g0 (.clr(clr), .Read1(w3), .Read2(w0), .Write(w10), .WriteData(WriteData), .clk(clk), .RegWrite(RegWrite), .Data1(rs), .Data2(rt));   //: @(390, 149) /sz:(147, 182) /sn:0 /p:[ Ti0>1 Li0>1 Li1>3 Li2>1 Li3>0 Bi0>1 Bi1>1 Ro0<1 Ro1<0 ]
  Extend g15 (.A(w8), .S(Inm32));   //: @(443, 447) /sz:(40, 40) /sn:0 /p:[ Li0>0 Ro0<0 ]
  //: input g13 (RegWrite) @(143,375) /sn:0 /w:[ 0 ]

endmodule

module Extend(S, A);
//: interface  /sz:(40, 40) /bd:[ Li0>A[15:0](23/40) Li1>A[15:0](23/40) Ro0<S[31:0](23/40) Ro1<S[31:0](23/40) ]
input [15:0] A;    //: /sn:0 {0}(307,243)(307,412)(325,412){1}
//: {2}(326,412)(355,412){3}
output [31:0] S;    //: /sn:0 /dp:1 {0}(361,332)(401,332){1}
wire w1;    //: /sn:0 {0}(326,407)(326,404){1}
//: {2}(328,402)(355,402){3}
//: {4}(326,400)(326,394){5}
//: {6}(328,392)(355,392){7}
//: {8}(326,390)(326,384){9}
//: {10}(328,382)(355,382){11}
//: {12}(326,380)(326,374){13}
//: {14}(328,372)(355,372){15}
//: {16}(326,370)(326,364){17}
//: {18}(328,362)(355,362){19}
//: {20}(326,360)(326,354){21}
//: {22}(328,352)(355,352){23}
//: {24}(326,350)(326,344){25}
//: {26}(328,342)(355,342){27}
//: {28}(326,340)(326,334){29}
//: {30}(328,332)(355,332){31}
//: {32}(326,330)(326,324){33}
//: {34}(328,322)(355,322){35}
//: {36}(326,320)(326,314){37}
//: {38}(328,312)(355,312){39}
//: {40}(326,310)(326,304){41}
//: {42}(328,302)(355,302){43}
//: {44}(326,300)(326,294){45}
//: {46}(328,292)(355,292){47}
//: {48}(326,290)(326,284){49}
//: {50}(328,282)(355,282){51}
//: {52}(326,280)(326,274){53}
//: {54}(328,272)(355,272){55}
//: {56}(326,270)(326,264){57}
//: {58}(328,262)(355,262){59}
//: {60}(326,260)(326,252)(355,252){61}
//: enddecls

  //: joint g8 (w1) @(326, 382) /w:[ 10 12 -1 9 ]
  tran g4(.Z(w1), .I(A[15]));   //: @(326,410) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:0
  //: joint g16 (w1) @(326, 302) /w:[ 42 44 -1 41 ]
  //: joint g17 (w1) @(326, 292) /w:[ 46 48 -1 45 ]
  concat g2 (.I0(A), .I1(w1), .I2(w1), .I3(w1), .I4(w1), .I5(w1), .I6(w1), .I7(w1), .I8(w1), .I9(w1), .I10(w1), .I11(w1), .I12(w1), .I13(w1), .I14(w1), .I15(w1), .I16(w1), .Z(S));   //: @(360,332) /sn:0 /w:[ 3 3 7 11 15 19 23 27 31 35 39 43 47 51 55 59 61 0 ] /dr:0
  //: output g1 (S) @(398,332) /sn:0 /w:[ 1 ]
  //: joint g18 (w1) @(326, 282) /w:[ 50 52 -1 49 ]
  //: joint g10 (w1) @(326, 362) /w:[ 18 20 -1 17 ]
  //: joint g9 (w1) @(326, 372) /w:[ 14 16 -1 13 ]
  //: joint g7 (w1) @(326, 392) /w:[ 6 8 -1 5 ]
  //: joint g12 (w1) @(326, 342) /w:[ 26 28 -1 25 ]
  //: joint g14 (w1) @(326, 322) /w:[ 34 36 -1 33 ]
  //: joint g11 (w1) @(326, 352) /w:[ 22 24 -1 21 ]
  //: joint g5 (w1) @(326, 402) /w:[ 2 4 -1 1 ]
  //: joint g19 (w1) @(326, 272) /w:[ 54 56 -1 53 ]
  //: joint g20 (w1) @(326, 262) /w:[ 58 60 -1 57 ]
  //: joint g15 (w1) @(326, 312) /w:[ 38 40 -1 37 ]
  //: input g0 (A) @(307,241) /sn:0 /R:3 /w:[ 0 ]
  //: joint g13 (w1) @(326, 332) /w:[ 30 32 -1 29 ]

endmodule

module main;    //: root_module
wire w13;    //: /sn:0 {0}(1365,410)(1365,137)(778,137){1}
wire [31:0] w6;    //: /sn:0 /dp:7 {0}(834,442)(728,442){1}
//: {2}(727,442)(724,442)(724,513){3}
//: {4}(724,514)(724,564)(711,564){5}
//: {6}(710,564)(687,564)(687,564)(680,564){7}
wire [31:0] w16;    //: /sn:0 /dp:1 {0}(1163,303)(1279,303)(1279,321)(1315,321){1}
wire [31:0] w7;    //: /sn:0 {0}(680,449)(692,449)(692,331)(1010,331){1}
//: {2}(1014,331)(1028,331){3}
//: {4}(1029,331)(1234,331){5}
//: {6}(1012,333)(1012,438)(1041,438){7}
wire Zero;    //: /sn:0 /dp:1 {0}(1185,444)(1213,444)(1213,246)(1248,246)(1248,256){1}
wire w25;    //: /sn:0 /dp:1 {0}(1851,264)(1851,324)(1750,324){1}
wire w4;    //: /sn:0 {0}(590,571)(523,571)(523,863){1}
//: {2}(525,865)(911,865)(911,632){3}
//: {4}(521,865)(483,865){5}
wire [31:0] Inm32;    //: /sn:0 /dp:1 {0}(973,561)(1041,561){1}
wire w22;    //: /sn:0 /dp:1 {0}(1811,217)(1811,290)(1750,290){1}
wire [5:0] w36;    //: /sn:0 {0}(1853,571)(1853,581)(1709,581)(1709,490){1}
wire w0;    //: /sn:0 {0}(1465,484)(1465,118)(778,118){1}
wire [31:0] w3;    //: /sn:0 /dp:1 {0}(1478,507)(1526,507)(1526,693)(868,693)(868,632){1}
wire w20;    //: /sn:0 {0}(778,69)(1331,69)(1331,308){1}
wire w29;    //: /sn:0 /dp:1 {0}(1889,312)(1889,359)(1750,359){1}
wire [25:0] w30;    //: /sn:0 {0}(711,559)(711,552)(774,552)(774,308)(1157,308){1}
wire [31:0] rt;    //: /sn:0 /dp:1 {0}(1041,527)(1018,527){1}
//: {2}(1014,527)(973,527){3}
//: {4}(1016,529)(1016,633)(1196,633)(1196,559)(1253,559){5}
wire w18;    //: /sn:0 /dp:1 {0}(1786,206)(1786,275)(1750,275){1}
wire w19;    //: /sn:0 {0}(778,84)(1253,84)(1253,256){1}
wire [31:0] w12;    //: /sn:0 {0}(1185,462)(1199,462)(1199,351)(1234,351){1}
wire [3:0] w23;    //: /sn:0 /dp:1 {0}(778,226)(1093,226)(1093,377)(1129,377)(1129,412){1}
wire w10;    //: /sn:0 /dp:1 {0}(1250,318)(1250,277){1}
wire [31:0] ALUResult;    //: /sn:0 /dp:1 {0}(1185,487)(1194,487)(1194,488)(1204,488){1}
//: {2}(1208,488)(1227,488){3}
//: {4}(1231,488)(1253,488){5}
//: {6}(1229,490)(1229,644)(1432,644)(1432,517)(1449,517){7}
//: {8}(1206,490)(1206,749)(1359,749)(1359,739){9}
wire w24;    //: /sn:0 /dp:1 {0}(1833,245)(1833,308)(1750,308){1}
wire w21;    //: /sn:0 {0}(1294,410)(1294,102)(778,102){1}
wire w31;    //: /sn:0 /dp:1 {0}(1903,334)(1903,378)(1750,378){1}
wire [31:0] w1;    //: /sn:0 {0}(1449,497)(1425,497)(1425,489)(1402,489){1}
wire RegDst;    //: /sn:0 {0}(834,533)(788,533)(788,261)(778,261){1}
wire w32;    //: /sn:0 /dp:1 {0}(1923,480)(1923,490)(1908,490)(1908,467)(1750,467){1}
wire w27;    //: /sn:0 {0}(778,172)(904,172)(904,411){1}
wire [5:0] w17;    //: /sn:0 {0}(728,514)(737,514)(737,284){1}
wire [3:0] w33;    //: /sn:0 /dp:1 {0}(1837,408)(1837,432)(1750,432){1}
wire w28;    //: /sn:0 /dp:1 {0}(1868,288)(1868,343)(1750,343){1}
wire [5:0] w35;    //: /sn:0 {0}(1606,563)(1606,573)(1682,573)(1682,490){1}
wire [31:0] w14;    //: /sn:0 /dp:1 {0}(1344,331)(1503,331)(1503,38)(582,38)(582,161){1}
//: {2}(580,163)(398,163)(398,101){3}
//: {4}(582,165)(582,424)(590,424){5}
wire [31:0] w11;    //: /sn:0 /dp:1 {0}(1263,341)(1315,341){1}
wire w2;    //: /sn:0 {0}(936,751)(936,632){1}
wire [5:0] w15;    //: /sn:0 {0}(1029,326)(1029,298)(1157,298){1}
wire [5:0] w5;    //: /sn:0 {0}(728,437)(728,430)(710,430)(710,284){1}
wire w26;    //: /sn:0 {0}(778,153)(1068,153)(1068,412){1}
wire w9;    //: /sn:0 {0}(522,455)(590,455){1}
wire [31:0] rs;    //: /sn:0 {0}(1041,494)(973,494){1}
//: enddecls

  //: joint g8 (w4) @(523, 865) /w:[ 2 1 4 -1 ]
  mux g4 (.I0(ALUResult), .I1(w1), .S(w0), .Z(w3));   //: @(1465,507) /sn:0 /R:1 /w:[ 7 0 0 0 ] /ss:1 /do:0
  Mem g3 (.MemRead(w21), .MemWrite(w13), .WriteData(rt), .Address(ALUResult), .ReadData(w1));   //: @(1254, 411) /sz:(147, 210) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>5 Li1>5 Ro0<1 ]
  tran g16(.Z(w15), .I(w7[31:26]));   //: @(1029,329) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:0
  //: dip g26 (w35) @(1606,553) /sn:0 /w:[ 0 ] /st:2
  //: comment g17 /dolink:0 /link:"" @(1319,280) /sn:0
  //: /line:"Jump"
  //: /end
  //: joint g2 (rt) @(1016, 527) /w:[ 1 -1 2 4 ]
  led g30 (.I(w24));   //: @(1833,238) /sn:0 /w:[ 0 ] /type:0
  tran g23(.Z(w17), .I(w6[5:0]));   //: @(722,514) /sn:0 /R:2 /w:[ 0 4 3 ] /ss:1
  and g24 (.I0(w19), .I1(Zero), .Z(w10));   //: @(1250,267) /sn:0 /R:3 /w:[ 1 1 1 ]
  EXE g1 (.ALUSrc(w26), .ALUOperation(w23), .PCNext(w7), .Inm32(Inm32), .rs(rs), .rt(rt), .BranchTarget(w12), .Zero(Zero), .ALUResult(ALUResult));   //: @(1042, 413) /sz:(142, 213) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>7 Li1>1 Li2>0 Li3>0 Ro0<0 Ro1<0 Ro2<0 ]
  led g39 (.I(ALUResult));   //: @(1359,732) /sn:0 /w:[ 9 ] /type:2
  led g29 (.I(w22));   //: @(1811,210) /sn:0 /w:[ 0 ] /type:0
  //: switch g18 (w2) @(936,765) /sn:0 /R:1 /w:[ 0 ] /st:1
  UC g25 (.Func(w36), .Op(w35), .RegDst(w32), .RegWrite(w31), .ALUSrc(w29), .MemWrite(w28), .ALUCtrl(w33), .MemToReg(w25), .MemRead(w24), .Jump(w18), .Branch(w22));   //: @(1648, 258) /sz:(101, 231) /sn:0 /p:[ Bi0>1 Bi1>1 Ro0<1 Ro1<1 Ro2<1 Ro3<1 Ro4<1 Ro5<1 Ro6<1 Ro7<1 Ro8<1 ]
  //: joint g10 (w7) @(1012, 331) /w:[ 2 -1 1 6 ]
  fetch g6 (.Reset(w9), .Clk(w4), .PCNew(w14), .PCNext(w7), .Inst(w6));   //: @(591, 411) /sz:(88, 222) /sn:0 /p:[ Li0>1 Li1>0 Li2>5 Ro0<0 Ro1<7 ]
  led g35 (.I(w32));   //: @(1923,473) /sn:0 /w:[ 0 ] /type:0
  clock g7 (.Z(w4));   //: @(470,865) /sn:0 /w:[ 5 ] /omega:6000 /phi:0 /duty:50
  led g31 (.I(w25));   //: @(1851,257) /sn:0 /w:[ 0 ] /type:0
  tran g22(.Z(w5), .I(w6[31:26]));   //: @(728,440) /sn:0 /R:1 /w:[ 0 2 1 ] /ss:0
  led g36 (.I(w33));   //: @(1837,401) /sn:0 /w:[ 0 ] /type:1
  led g33 (.I(w29));   //: @(1889,305) /sn:0 /w:[ 0 ] /type:0
  //: joint g40 (ALUResult) @(1206, 488) /w:[ 2 -1 1 8 ]
  //: comment g12 /dolink:0 /link:"" @(1219,282) /sn:0
  //: /line:"PCSrc"
  //: /end
  led g34 (.I(w31));   //: @(1903,327) /sn:0 /w:[ 0 ] /type:0
  led g28 (.I(w18));   //: @(1786,199) /sn:0 /w:[ 0 ] /type:0
  //: joint g5 (ALUResult) @(1229, 488) /w:[ 4 -1 3 6 ]
  mux g11 (.I0(w7), .I1(w12), .S(w10), .Z(w11));   //: @(1250,341) /sn:0 /R:1 /w:[ 5 1 0 0 ] /ss:1 /do:1
  concat g14 (.I0(w30), .I1(w15), .Z(w16));   //: @(1162,303) /sn:0 /w:[ 1 1 0 ] /dr:0
  UC g21 (.Func(w17), .Op(w5), .RegDst(RegDst), .RegWrite(w27), .ALUSrc(w26), .MemWrite(w13), .ALUCtrl(w23), .MemToReg(w0), .MemRead(w21), .Jump(w20), .Branch(w19));   //: @(676, 52) /sz:(101, 231) /sn:0 /p:[ Bi0>1 Bi1>1 Ro0<1 Ro1<0 Ro2<0 Ro3<1 Ro4<0 Ro5<1 Ro6<1 Ro7<0 Ro8<0 ]
  //: switch g19 (w9) @(505,455) /sn:0 /w:[ 0 ] /st:0
  led g32 (.I(w28));   //: @(1868,281) /sn:0 /w:[ 0 ] /type:0
  //: comment g20 /dolink:0 /link:"" @(1473,465) /sn:0
  //: /line:"MemtoReg"
  //: /end
  Read g0 (.RegWrite(w27), .RegDst(RegDst), .Inst(w6), .clk(w4), .clr(w2), .WriteData(w3), .Inm32(Inm32), .rt(rt), .rs(rs));   //: @(835, 412) /sz:(137, 219) /sn:0 /p:[ Ti0>1 Li0>0 Li1>0 Bi0>3 Bi1>1 Bi2>1 Ro0<0 Ro1<3 Ro2<1 ]
  //: joint g38 (w14) @(582, 163) /w:[ -1 1 2 4 ]
  tran g15(.Z(w30), .I(w6[25:0]));   //: @(711,562) /sn:0 /R:1 /w:[ 0 6 5 ] /ss:0
  //: dip g27 (w36) @(1853,561) /sn:0 /w:[ 0 ] /st:0
  led g37 (.I(w14));   //: @(398,94) /sn:0 /w:[ 3 ] /type:2
  mux g13 (.I0(w11), .I1(w16), .S(w20), .Z(w14));   //: @(1331,331) /sn:0 /R:1 /w:[ 1 1 1 0 ] /ss:1 /do:0

endmodule
